module LookupTable(
  input         clock,
  input         reset,
  output [31:0] io_data_0,
  output [31:0] io_data_1,
  output [31:0] io_data_2,
  output [31:0] io_data_3,
  output [31:0] io_data_4,
  output [31:0] io_data_5,
  output [31:0] io_data_6,
  output [31:0] io_data_7,
  output [31:0] io_data_8,
  output [31:0] io_data_9,
  output [31:0] io_data_10,
  output [31:0] io_data_11,
  output [31:0] io_data_12,
  output [31:0] io_data_13,
  input  [31:0] io_dataIn_0,
  input  [31:0] io_dataIn_1,
  input         io_writeFlag_0,
  input         io_writeFlag_1,
  input  [4:0]  io_wptr_0,
  input  [4:0]  io_wptr_1,
  input  [63:0] config_awaddr,
  input         config_awvalid,
  output        config_awready,
  input  [63:0] config_araddr,
  input         config_arvalid,
  output        config_arready,
  input  [31:0] config_wdata,
  input         config_wvalid,
  output        config_wready,
  output [31:0] config_rdata,
  output        config_rvalid,
  input         config_rready,
  output        config_bvalid,
  input         config_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] table_0; // @[util.scala 16:22]
  reg [31:0] table_1; // @[util.scala 16:22]
  reg [31:0] table_2; // @[util.scala 16:22]
  reg [31:0] table_3; // @[util.scala 16:22]
  reg [31:0] table_4; // @[util.scala 16:22]
  reg [31:0] table_5; // @[util.scala 16:22]
  reg [31:0] table_6; // @[util.scala 16:22]
  reg [31:0] table_7; // @[util.scala 16:22]
  reg [31:0] table_8; // @[util.scala 16:22]
  reg [31:0] table_9; // @[util.scala 16:22]
  reg [31:0] table_10; // @[util.scala 16:22]
  reg [31:0] table_11; // @[util.scala 16:22]
  reg [31:0] table_12; // @[util.scala 16:22]
  reg [31:0] table_13; // @[util.scala 16:22]
  reg [31:0] table_14; // @[util.scala 16:22]
  reg [31:0] table_15; // @[util.scala 16:22]
  reg [31:0] table_16; // @[util.scala 16:22]
  reg [31:0] table_17; // @[util.scala 16:22]
  reg [31:0] table_18; // @[util.scala 16:22]
  reg [31:0] table_19; // @[util.scala 16:22]
  reg [31:0] table_20; // @[util.scala 16:22]
  reg [31:0] table_21; // @[util.scala 16:22]
  reg [31:0] table_22; // @[util.scala 16:22]
  reg [31:0] table_23; // @[util.scala 16:22]
  reg [31:0] table_24; // @[util.scala 16:22]
  reg [31:0] table_25; // @[util.scala 16:22]
  reg [31:0] table_26; // @[util.scala 16:22]
  reg [31:0] table_27; // @[util.scala 16:22]
  reg [31:0] table_28; // @[util.scala 16:22]
  reg [31:0] table_29; // @[util.scala 16:22]
  reg [31:0] table_30; // @[util.scala 16:22]
  reg [31:0] table_31; // @[util.scala 16:22]
  reg [2:0] status; // @[util.scala 26:23]
  wire [2:0] _GEN_3 = config_bready ? 3'h0 : status; // @[util.scala 41:24 util.scala 42:14 util.scala 26:23]
  wire [2:0] _GEN_4 = config_rready ? 3'h0 : status; // @[util.scala 47:25 util.scala 48:14 util.scala 26:23]
  wire [2:0] _GEN_5 = status == 3'h5 ? _GEN_4 : status; // @[util.scala 46:36 util.scala 26:23]
  wire [2:0] _GEN_6 = status == 3'h4 ? 3'h5 : _GEN_5; // @[util.scala 44:35 util.scala 45:12]
  wire [2:0] _GEN_7 = status == 3'h3 ? _GEN_3 : _GEN_6; // @[util.scala 40:35]
  wire  wvalid = config_wvalid & config_wready; // @[util.scala 64:30]
  reg [4:0] ewaddr; // @[util.scala 65:19]
  wire  _T_7 = io_writeFlag_0 & io_writeFlag_1; // @[util.scala 70:39]
  wire [31:0] _GEN_12 = 5'h0 == ewaddr ? config_wdata : table_0; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_13 = 5'h1 == ewaddr ? config_wdata : table_1; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_14 = 5'h2 == ewaddr ? config_wdata : table_2; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_15 = 5'h3 == ewaddr ? config_wdata : table_3; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_16 = 5'h4 == ewaddr ? config_wdata : table_4; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_17 = 5'h5 == ewaddr ? config_wdata : table_5; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_18 = 5'h6 == ewaddr ? config_wdata : table_6; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_19 = 5'h7 == ewaddr ? config_wdata : table_7; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_20 = 5'h8 == ewaddr ? config_wdata : table_8; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_21 = 5'h9 == ewaddr ? config_wdata : table_9; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_22 = 5'ha == ewaddr ? config_wdata : table_10; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_23 = 5'hb == ewaddr ? config_wdata : table_11; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_24 = 5'hc == ewaddr ? config_wdata : table_12; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_25 = 5'hd == ewaddr ? config_wdata : table_13; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_26 = 5'he == ewaddr ? config_wdata : table_14; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_27 = 5'hf == ewaddr ? config_wdata : table_15; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_28 = 5'h10 == ewaddr ? config_wdata : table_16; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_29 = 5'h11 == ewaddr ? config_wdata : table_17; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_30 = 5'h12 == ewaddr ? config_wdata : table_18; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_31 = 5'h13 == ewaddr ? config_wdata : table_19; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_32 = 5'h14 == ewaddr ? config_wdata : table_20; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_33 = 5'h15 == ewaddr ? config_wdata : table_21; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_34 = 5'h16 == ewaddr ? config_wdata : table_22; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_35 = 5'h17 == ewaddr ? config_wdata : table_23; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_36 = 5'h18 == ewaddr ? config_wdata : table_24; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_37 = 5'h19 == ewaddr ? config_wdata : table_25; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_38 = 5'h1a == ewaddr ? config_wdata : table_26; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_39 = 5'h1b == ewaddr ? config_wdata : table_27; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_40 = 5'h1c == ewaddr ? config_wdata : table_28; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_41 = 5'h1d == ewaddr ? config_wdata : table_29; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_42 = 5'h1e == ewaddr ? config_wdata : table_30; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_43 = 5'h1f == ewaddr ? config_wdata : table_31; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_44 = 5'h0 == io_wptr_0 ? io_dataIn_0 : _GEN_12; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_45 = 5'h1 == io_wptr_0 ? io_dataIn_0 : _GEN_13; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_46 = 5'h2 == io_wptr_0 ? io_dataIn_0 : _GEN_14; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_47 = 5'h3 == io_wptr_0 ? io_dataIn_0 : _GEN_15; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_48 = 5'h4 == io_wptr_0 ? io_dataIn_0 : _GEN_16; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_49 = 5'h5 == io_wptr_0 ? io_dataIn_0 : _GEN_17; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_50 = 5'h6 == io_wptr_0 ? io_dataIn_0 : _GEN_18; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_51 = 5'h7 == io_wptr_0 ? io_dataIn_0 : _GEN_19; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_52 = 5'h8 == io_wptr_0 ? io_dataIn_0 : _GEN_20; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_53 = 5'h9 == io_wptr_0 ? io_dataIn_0 : _GEN_21; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_54 = 5'ha == io_wptr_0 ? io_dataIn_0 : _GEN_22; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_55 = 5'hb == io_wptr_0 ? io_dataIn_0 : _GEN_23; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_56 = 5'hc == io_wptr_0 ? io_dataIn_0 : _GEN_24; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_57 = 5'hd == io_wptr_0 ? io_dataIn_0 : _GEN_25; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_58 = 5'he == io_wptr_0 ? io_dataIn_0 : _GEN_26; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_59 = 5'hf == io_wptr_0 ? io_dataIn_0 : _GEN_27; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_60 = 5'h10 == io_wptr_0 ? io_dataIn_0 : _GEN_28; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_61 = 5'h11 == io_wptr_0 ? io_dataIn_0 : _GEN_29; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_62 = 5'h12 == io_wptr_0 ? io_dataIn_0 : _GEN_30; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_63 = 5'h13 == io_wptr_0 ? io_dataIn_0 : _GEN_31; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_64 = 5'h14 == io_wptr_0 ? io_dataIn_0 : _GEN_32; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_65 = 5'h15 == io_wptr_0 ? io_dataIn_0 : _GEN_33; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_66 = 5'h16 == io_wptr_0 ? io_dataIn_0 : _GEN_34; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_67 = 5'h17 == io_wptr_0 ? io_dataIn_0 : _GEN_35; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_68 = 5'h18 == io_wptr_0 ? io_dataIn_0 : _GEN_36; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_69 = 5'h19 == io_wptr_0 ? io_dataIn_0 : _GEN_37; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_70 = 5'h1a == io_wptr_0 ? io_dataIn_0 : _GEN_38; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_71 = 5'h1b == io_wptr_0 ? io_dataIn_0 : _GEN_39; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_72 = 5'h1c == io_wptr_0 ? io_dataIn_0 : _GEN_40; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_73 = 5'h1d == io_wptr_0 ? io_dataIn_0 : _GEN_41; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_74 = 5'h1e == io_wptr_0 ? io_dataIn_0 : _GEN_42; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_75 = 5'h1f == io_wptr_0 ? io_dataIn_0 : _GEN_43; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_204 = 5'h0 == io_wptr_1 ? io_dataIn_1 : _GEN_12; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_205 = 5'h1 == io_wptr_1 ? io_dataIn_1 : _GEN_13; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_206 = 5'h2 == io_wptr_1 ? io_dataIn_1 : _GEN_14; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_207 = 5'h3 == io_wptr_1 ? io_dataIn_1 : _GEN_15; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_208 = 5'h4 == io_wptr_1 ? io_dataIn_1 : _GEN_16; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_209 = 5'h5 == io_wptr_1 ? io_dataIn_1 : _GEN_17; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_210 = 5'h6 == io_wptr_1 ? io_dataIn_1 : _GEN_18; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_211 = 5'h7 == io_wptr_1 ? io_dataIn_1 : _GEN_19; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_212 = 5'h8 == io_wptr_1 ? io_dataIn_1 : _GEN_20; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_213 = 5'h9 == io_wptr_1 ? io_dataIn_1 : _GEN_21; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_214 = 5'ha == io_wptr_1 ? io_dataIn_1 : _GEN_22; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_215 = 5'hb == io_wptr_1 ? io_dataIn_1 : _GEN_23; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_216 = 5'hc == io_wptr_1 ? io_dataIn_1 : _GEN_24; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_217 = 5'hd == io_wptr_1 ? io_dataIn_1 : _GEN_25; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_218 = 5'he == io_wptr_1 ? io_dataIn_1 : _GEN_26; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_219 = 5'hf == io_wptr_1 ? io_dataIn_1 : _GEN_27; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_220 = 5'h10 == io_wptr_1 ? io_dataIn_1 : _GEN_28; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_221 = 5'h11 == io_wptr_1 ? io_dataIn_1 : _GEN_29; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_222 = 5'h12 == io_wptr_1 ? io_dataIn_1 : _GEN_30; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_223 = 5'h13 == io_wptr_1 ? io_dataIn_1 : _GEN_31; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_224 = 5'h14 == io_wptr_1 ? io_dataIn_1 : _GEN_32; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_225 = 5'h15 == io_wptr_1 ? io_dataIn_1 : _GEN_33; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_226 = 5'h16 == io_wptr_1 ? io_dataIn_1 : _GEN_34; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_227 = 5'h17 == io_wptr_1 ? io_dataIn_1 : _GEN_35; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_228 = 5'h18 == io_wptr_1 ? io_dataIn_1 : _GEN_36; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_229 = 5'h19 == io_wptr_1 ? io_dataIn_1 : _GEN_37; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_230 = 5'h1a == io_wptr_1 ? io_dataIn_1 : _GEN_38; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_231 = 5'h1b == io_wptr_1 ? io_dataIn_1 : _GEN_39; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_232 = 5'h1c == io_wptr_1 ? io_dataIn_1 : _GEN_40; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_233 = 5'h1d == io_wptr_1 ? io_dataIn_1 : _GEN_41; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_234 = 5'h1e == io_wptr_1 ? io_dataIn_1 : _GEN_42; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_235 = 5'h1f == io_wptr_1 ? io_dataIn_1 : _GEN_43; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_268 = 5'h0 == io_wptr_0 ? io_dataIn_0 : table_0; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_269 = 5'h1 == io_wptr_0 ? io_dataIn_0 : table_1; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_270 = 5'h2 == io_wptr_0 ? io_dataIn_0 : table_2; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_271 = 5'h3 == io_wptr_0 ? io_dataIn_0 : table_3; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_272 = 5'h4 == io_wptr_0 ? io_dataIn_0 : table_4; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_273 = 5'h5 == io_wptr_0 ? io_dataIn_0 : table_5; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_274 = 5'h6 == io_wptr_0 ? io_dataIn_0 : table_6; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_275 = 5'h7 == io_wptr_0 ? io_dataIn_0 : table_7; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_276 = 5'h8 == io_wptr_0 ? io_dataIn_0 : table_8; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_277 = 5'h9 == io_wptr_0 ? io_dataIn_0 : table_9; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_278 = 5'ha == io_wptr_0 ? io_dataIn_0 : table_10; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_279 = 5'hb == io_wptr_0 ? io_dataIn_0 : table_11; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_280 = 5'hc == io_wptr_0 ? io_dataIn_0 : table_12; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_281 = 5'hd == io_wptr_0 ? io_dataIn_0 : table_13; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_282 = 5'he == io_wptr_0 ? io_dataIn_0 : table_14; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_283 = 5'hf == io_wptr_0 ? io_dataIn_0 : table_15; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_284 = 5'h10 == io_wptr_0 ? io_dataIn_0 : table_16; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_285 = 5'h11 == io_wptr_0 ? io_dataIn_0 : table_17; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_286 = 5'h12 == io_wptr_0 ? io_dataIn_0 : table_18; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_287 = 5'h13 == io_wptr_0 ? io_dataIn_0 : table_19; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_288 = 5'h14 == io_wptr_0 ? io_dataIn_0 : table_20; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_289 = 5'h15 == io_wptr_0 ? io_dataIn_0 : table_21; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_290 = 5'h16 == io_wptr_0 ? io_dataIn_0 : table_22; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_291 = 5'h17 == io_wptr_0 ? io_dataIn_0 : table_23; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_292 = 5'h18 == io_wptr_0 ? io_dataIn_0 : table_24; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_293 = 5'h19 == io_wptr_0 ? io_dataIn_0 : table_25; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_294 = 5'h1a == io_wptr_0 ? io_dataIn_0 : table_26; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_295 = 5'h1b == io_wptr_0 ? io_dataIn_0 : table_27; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_296 = 5'h1c == io_wptr_0 ? io_dataIn_0 : table_28; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_297 = 5'h1d == io_wptr_0 ? io_dataIn_0 : table_29; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_298 = 5'h1e == io_wptr_0 ? io_dataIn_0 : table_30; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_299 = 5'h1f == io_wptr_0 ? io_dataIn_0 : table_31; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_300 = 5'h0 == io_wptr_1 ? io_dataIn_1 : _GEN_268; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_301 = 5'h1 == io_wptr_1 ? io_dataIn_1 : _GEN_269; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_302 = 5'h2 == io_wptr_1 ? io_dataIn_1 : _GEN_270; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_303 = 5'h3 == io_wptr_1 ? io_dataIn_1 : _GEN_271; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_304 = 5'h4 == io_wptr_1 ? io_dataIn_1 : _GEN_272; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_305 = 5'h5 == io_wptr_1 ? io_dataIn_1 : _GEN_273; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_306 = 5'h6 == io_wptr_1 ? io_dataIn_1 : _GEN_274; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_307 = 5'h7 == io_wptr_1 ? io_dataIn_1 : _GEN_275; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_308 = 5'h8 == io_wptr_1 ? io_dataIn_1 : _GEN_276; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_309 = 5'h9 == io_wptr_1 ? io_dataIn_1 : _GEN_277; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_310 = 5'ha == io_wptr_1 ? io_dataIn_1 : _GEN_278; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_311 = 5'hb == io_wptr_1 ? io_dataIn_1 : _GEN_279; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_312 = 5'hc == io_wptr_1 ? io_dataIn_1 : _GEN_280; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_313 = 5'hd == io_wptr_1 ? io_dataIn_1 : _GEN_281; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_314 = 5'he == io_wptr_1 ? io_dataIn_1 : _GEN_282; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_315 = 5'hf == io_wptr_1 ? io_dataIn_1 : _GEN_283; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_316 = 5'h10 == io_wptr_1 ? io_dataIn_1 : _GEN_284; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_317 = 5'h11 == io_wptr_1 ? io_dataIn_1 : _GEN_285; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_318 = 5'h12 == io_wptr_1 ? io_dataIn_1 : _GEN_286; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_319 = 5'h13 == io_wptr_1 ? io_dataIn_1 : _GEN_287; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_320 = 5'h14 == io_wptr_1 ? io_dataIn_1 : _GEN_288; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_321 = 5'h15 == io_wptr_1 ? io_dataIn_1 : _GEN_289; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_322 = 5'h16 == io_wptr_1 ? io_dataIn_1 : _GEN_290; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_323 = 5'h17 == io_wptr_1 ? io_dataIn_1 : _GEN_291; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_324 = 5'h18 == io_wptr_1 ? io_dataIn_1 : _GEN_292; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_325 = 5'h19 == io_wptr_1 ? io_dataIn_1 : _GEN_293; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_326 = 5'h1a == io_wptr_1 ? io_dataIn_1 : _GEN_294; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_327 = 5'h1b == io_wptr_1 ? io_dataIn_1 : _GEN_295; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_328 = 5'h1c == io_wptr_1 ? io_dataIn_1 : _GEN_296; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_329 = 5'h1d == io_wptr_1 ? io_dataIn_1 : _GEN_297; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_330 = 5'h1e == io_wptr_1 ? io_dataIn_1 : _GEN_298; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_331 = 5'h1f == io_wptr_1 ? io_dataIn_1 : _GEN_299; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_364 = 5'h0 == io_wptr_1 ? io_dataIn_1 : table_0; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_365 = 5'h1 == io_wptr_1 ? io_dataIn_1 : table_1; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_366 = 5'h2 == io_wptr_1 ? io_dataIn_1 : table_2; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_367 = 5'h3 == io_wptr_1 ? io_dataIn_1 : table_3; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_368 = 5'h4 == io_wptr_1 ? io_dataIn_1 : table_4; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_369 = 5'h5 == io_wptr_1 ? io_dataIn_1 : table_5; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_370 = 5'h6 == io_wptr_1 ? io_dataIn_1 : table_6; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_371 = 5'h7 == io_wptr_1 ? io_dataIn_1 : table_7; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_372 = 5'h8 == io_wptr_1 ? io_dataIn_1 : table_8; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_373 = 5'h9 == io_wptr_1 ? io_dataIn_1 : table_9; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_374 = 5'ha == io_wptr_1 ? io_dataIn_1 : table_10; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_375 = 5'hb == io_wptr_1 ? io_dataIn_1 : table_11; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_376 = 5'hc == io_wptr_1 ? io_dataIn_1 : table_12; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_377 = 5'hd == io_wptr_1 ? io_dataIn_1 : table_13; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_378 = 5'he == io_wptr_1 ? io_dataIn_1 : table_14; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_379 = 5'hf == io_wptr_1 ? io_dataIn_1 : table_15; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_380 = 5'h10 == io_wptr_1 ? io_dataIn_1 : table_16; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_381 = 5'h11 == io_wptr_1 ? io_dataIn_1 : table_17; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_382 = 5'h12 == io_wptr_1 ? io_dataIn_1 : table_18; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_383 = 5'h13 == io_wptr_1 ? io_dataIn_1 : table_19; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_384 = 5'h14 == io_wptr_1 ? io_dataIn_1 : table_20; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_385 = 5'h15 == io_wptr_1 ? io_dataIn_1 : table_21; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_386 = 5'h16 == io_wptr_1 ? io_dataIn_1 : table_22; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_387 = 5'h17 == io_wptr_1 ? io_dataIn_1 : table_23; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_388 = 5'h18 == io_wptr_1 ? io_dataIn_1 : table_24; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_389 = 5'h19 == io_wptr_1 ? io_dataIn_1 : table_25; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_390 = 5'h1a == io_wptr_1 ? io_dataIn_1 : table_26; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_391 = 5'h1b == io_wptr_1 ? io_dataIn_1 : table_27; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_392 = 5'h1c == io_wptr_1 ? io_dataIn_1 : table_28; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_393 = 5'h1d == io_wptr_1 ? io_dataIn_1 : table_29; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_394 = 5'h1e == io_wptr_1 ? io_dataIn_1 : table_30; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_395 = 5'h1f == io_wptr_1 ? io_dataIn_1 : table_31; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_396 = io_writeFlag_1 ? _GEN_364 : table_0; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_397 = io_writeFlag_1 ? _GEN_365 : table_1; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_398 = io_writeFlag_1 ? _GEN_366 : table_2; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_399 = io_writeFlag_1 ? _GEN_367 : table_3; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_400 = io_writeFlag_1 ? _GEN_368 : table_4; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_401 = io_writeFlag_1 ? _GEN_369 : table_5; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_402 = io_writeFlag_1 ? _GEN_370 : table_6; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_403 = io_writeFlag_1 ? _GEN_371 : table_7; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_404 = io_writeFlag_1 ? _GEN_372 : table_8; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_405 = io_writeFlag_1 ? _GEN_373 : table_9; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_406 = io_writeFlag_1 ? _GEN_374 : table_10; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_407 = io_writeFlag_1 ? _GEN_375 : table_11; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_408 = io_writeFlag_1 ? _GEN_376 : table_12; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_409 = io_writeFlag_1 ? _GEN_377 : table_13; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_410 = io_writeFlag_1 ? _GEN_378 : table_14; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_411 = io_writeFlag_1 ? _GEN_379 : table_15; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_412 = io_writeFlag_1 ? _GEN_380 : table_16; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_413 = io_writeFlag_1 ? _GEN_381 : table_17; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_414 = io_writeFlag_1 ? _GEN_382 : table_18; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_415 = io_writeFlag_1 ? _GEN_383 : table_19; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_416 = io_writeFlag_1 ? _GEN_384 : table_20; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_417 = io_writeFlag_1 ? _GEN_385 : table_21; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_418 = io_writeFlag_1 ? _GEN_386 : table_22; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_419 = io_writeFlag_1 ? _GEN_387 : table_23; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_420 = io_writeFlag_1 ? _GEN_388 : table_24; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_421 = io_writeFlag_1 ? _GEN_389 : table_25; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_422 = io_writeFlag_1 ? _GEN_390 : table_26; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_423 = io_writeFlag_1 ? _GEN_391 : table_27; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_424 = io_writeFlag_1 ? _GEN_392 : table_28; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_425 = io_writeFlag_1 ? _GEN_393 : table_29; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_426 = io_writeFlag_1 ? _GEN_394 : table_30; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_427 = io_writeFlag_1 ? _GEN_395 : table_31; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_428 = io_writeFlag_0 ? _GEN_268 : _GEN_396; // @[util.scala 85:30]
  wire [31:0] _GEN_429 = io_writeFlag_0 ? _GEN_269 : _GEN_397; // @[util.scala 85:30]
  wire [31:0] _GEN_430 = io_writeFlag_0 ? _GEN_270 : _GEN_398; // @[util.scala 85:30]
  wire [31:0] _GEN_431 = io_writeFlag_0 ? _GEN_271 : _GEN_399; // @[util.scala 85:30]
  wire [31:0] _GEN_432 = io_writeFlag_0 ? _GEN_272 : _GEN_400; // @[util.scala 85:30]
  wire [31:0] _GEN_433 = io_writeFlag_0 ? _GEN_273 : _GEN_401; // @[util.scala 85:30]
  wire [31:0] _GEN_434 = io_writeFlag_0 ? _GEN_274 : _GEN_402; // @[util.scala 85:30]
  wire [31:0] _GEN_435 = io_writeFlag_0 ? _GEN_275 : _GEN_403; // @[util.scala 85:30]
  wire [31:0] _GEN_436 = io_writeFlag_0 ? _GEN_276 : _GEN_404; // @[util.scala 85:30]
  wire [31:0] _GEN_437 = io_writeFlag_0 ? _GEN_277 : _GEN_405; // @[util.scala 85:30]
  wire [31:0] _GEN_438 = io_writeFlag_0 ? _GEN_278 : _GEN_406; // @[util.scala 85:30]
  wire [31:0] _GEN_439 = io_writeFlag_0 ? _GEN_279 : _GEN_407; // @[util.scala 85:30]
  wire [31:0] _GEN_440 = io_writeFlag_0 ? _GEN_280 : _GEN_408; // @[util.scala 85:30]
  wire [31:0] _GEN_441 = io_writeFlag_0 ? _GEN_281 : _GEN_409; // @[util.scala 85:30]
  wire [31:0] _GEN_442 = io_writeFlag_0 ? _GEN_282 : _GEN_410; // @[util.scala 85:30]
  wire [31:0] _GEN_443 = io_writeFlag_0 ? _GEN_283 : _GEN_411; // @[util.scala 85:30]
  wire [31:0] _GEN_444 = io_writeFlag_0 ? _GEN_284 : _GEN_412; // @[util.scala 85:30]
  wire [31:0] _GEN_445 = io_writeFlag_0 ? _GEN_285 : _GEN_413; // @[util.scala 85:30]
  wire [31:0] _GEN_446 = io_writeFlag_0 ? _GEN_286 : _GEN_414; // @[util.scala 85:30]
  wire [31:0] _GEN_447 = io_writeFlag_0 ? _GEN_287 : _GEN_415; // @[util.scala 85:30]
  wire [31:0] _GEN_448 = io_writeFlag_0 ? _GEN_288 : _GEN_416; // @[util.scala 85:30]
  wire [31:0] _GEN_449 = io_writeFlag_0 ? _GEN_289 : _GEN_417; // @[util.scala 85:30]
  wire [31:0] _GEN_450 = io_writeFlag_0 ? _GEN_290 : _GEN_418; // @[util.scala 85:30]
  wire [31:0] _GEN_451 = io_writeFlag_0 ? _GEN_291 : _GEN_419; // @[util.scala 85:30]
  wire [31:0] _GEN_452 = io_writeFlag_0 ? _GEN_292 : _GEN_420; // @[util.scala 85:30]
  wire [31:0] _GEN_453 = io_writeFlag_0 ? _GEN_293 : _GEN_421; // @[util.scala 85:30]
  wire [31:0] _GEN_454 = io_writeFlag_0 ? _GEN_294 : _GEN_422; // @[util.scala 85:30]
  wire [31:0] _GEN_455 = io_writeFlag_0 ? _GEN_295 : _GEN_423; // @[util.scala 85:30]
  wire [31:0] _GEN_456 = io_writeFlag_0 ? _GEN_296 : _GEN_424; // @[util.scala 85:30]
  wire [31:0] _GEN_457 = io_writeFlag_0 ? _GEN_297 : _GEN_425; // @[util.scala 85:30]
  wire [31:0] _GEN_458 = io_writeFlag_0 ? _GEN_298 : _GEN_426; // @[util.scala 85:30]
  wire [31:0] _GEN_459 = io_writeFlag_0 ? _GEN_299 : _GEN_427; // @[util.scala 85:30]
  wire [31:0] _GEN_460 = _T_7 ? _GEN_300 : _GEN_428; // @[util.scala 82:39]
  wire [31:0] _GEN_461 = _T_7 ? _GEN_301 : _GEN_429; // @[util.scala 82:39]
  wire [31:0] _GEN_462 = _T_7 ? _GEN_302 : _GEN_430; // @[util.scala 82:39]
  wire [31:0] _GEN_463 = _T_7 ? _GEN_303 : _GEN_431; // @[util.scala 82:39]
  wire [31:0] _GEN_464 = _T_7 ? _GEN_304 : _GEN_432; // @[util.scala 82:39]
  wire [31:0] _GEN_465 = _T_7 ? _GEN_305 : _GEN_433; // @[util.scala 82:39]
  wire [31:0] _GEN_466 = _T_7 ? _GEN_306 : _GEN_434; // @[util.scala 82:39]
  wire [31:0] _GEN_467 = _T_7 ? _GEN_307 : _GEN_435; // @[util.scala 82:39]
  wire [31:0] _GEN_468 = _T_7 ? _GEN_308 : _GEN_436; // @[util.scala 82:39]
  wire [31:0] _GEN_469 = _T_7 ? _GEN_309 : _GEN_437; // @[util.scala 82:39]
  wire [31:0] _GEN_470 = _T_7 ? _GEN_310 : _GEN_438; // @[util.scala 82:39]
  wire [31:0] _GEN_471 = _T_7 ? _GEN_311 : _GEN_439; // @[util.scala 82:39]
  wire [31:0] _GEN_472 = _T_7 ? _GEN_312 : _GEN_440; // @[util.scala 82:39]
  wire [31:0] _GEN_473 = _T_7 ? _GEN_313 : _GEN_441; // @[util.scala 82:39]
  wire [31:0] _GEN_474 = _T_7 ? _GEN_314 : _GEN_442; // @[util.scala 82:39]
  wire [31:0] _GEN_475 = _T_7 ? _GEN_315 : _GEN_443; // @[util.scala 82:39]
  wire [31:0] _GEN_476 = _T_7 ? _GEN_316 : _GEN_444; // @[util.scala 82:39]
  wire [31:0] _GEN_477 = _T_7 ? _GEN_317 : _GEN_445; // @[util.scala 82:39]
  wire [31:0] _GEN_478 = _T_7 ? _GEN_318 : _GEN_446; // @[util.scala 82:39]
  wire [31:0] _GEN_479 = _T_7 ? _GEN_319 : _GEN_447; // @[util.scala 82:39]
  wire [31:0] _GEN_480 = _T_7 ? _GEN_320 : _GEN_448; // @[util.scala 82:39]
  wire [31:0] _GEN_481 = _T_7 ? _GEN_321 : _GEN_449; // @[util.scala 82:39]
  wire [31:0] _GEN_482 = _T_7 ? _GEN_322 : _GEN_450; // @[util.scala 82:39]
  wire [31:0] _GEN_483 = _T_7 ? _GEN_323 : _GEN_451; // @[util.scala 82:39]
  wire [31:0] _GEN_484 = _T_7 ? _GEN_324 : _GEN_452; // @[util.scala 82:39]
  wire [31:0] _GEN_485 = _T_7 ? _GEN_325 : _GEN_453; // @[util.scala 82:39]
  wire [31:0] _GEN_486 = _T_7 ? _GEN_326 : _GEN_454; // @[util.scala 82:39]
  wire [31:0] _GEN_487 = _T_7 ? _GEN_327 : _GEN_455; // @[util.scala 82:39]
  wire [31:0] _GEN_488 = _T_7 ? _GEN_328 : _GEN_456; // @[util.scala 82:39]
  wire [31:0] _GEN_489 = _T_7 ? _GEN_329 : _GEN_457; // @[util.scala 82:39]
  wire [31:0] _GEN_490 = _T_7 ? _GEN_330 : _GEN_458; // @[util.scala 82:39]
  wire [31:0] _GEN_491 = _T_7 ? _GEN_331 : _GEN_459; // @[util.scala 82:39]
  wire [31:0] _GEN_492 = wvalid ? _GEN_12 : _GEN_460; // @[util.scala 80:21]
  wire [31:0] _GEN_493 = wvalid ? _GEN_13 : _GEN_461; // @[util.scala 80:21]
  wire [31:0] _GEN_494 = wvalid ? _GEN_14 : _GEN_462; // @[util.scala 80:21]
  wire [31:0] _GEN_495 = wvalid ? _GEN_15 : _GEN_463; // @[util.scala 80:21]
  wire [31:0] _GEN_496 = wvalid ? _GEN_16 : _GEN_464; // @[util.scala 80:21]
  wire [31:0] _GEN_497 = wvalid ? _GEN_17 : _GEN_465; // @[util.scala 80:21]
  wire [31:0] _GEN_498 = wvalid ? _GEN_18 : _GEN_466; // @[util.scala 80:21]
  wire [31:0] _GEN_499 = wvalid ? _GEN_19 : _GEN_467; // @[util.scala 80:21]
  wire [31:0] _GEN_500 = wvalid ? _GEN_20 : _GEN_468; // @[util.scala 80:21]
  wire [31:0] _GEN_501 = wvalid ? _GEN_21 : _GEN_469; // @[util.scala 80:21]
  wire [31:0] _GEN_502 = wvalid ? _GEN_22 : _GEN_470; // @[util.scala 80:21]
  wire [31:0] _GEN_503 = wvalid ? _GEN_23 : _GEN_471; // @[util.scala 80:21]
  wire [31:0] _GEN_504 = wvalid ? _GEN_24 : _GEN_472; // @[util.scala 80:21]
  wire [31:0] _GEN_505 = wvalid ? _GEN_25 : _GEN_473; // @[util.scala 80:21]
  wire [31:0] _GEN_506 = wvalid ? _GEN_26 : _GEN_474; // @[util.scala 80:21]
  wire [31:0] _GEN_507 = wvalid ? _GEN_27 : _GEN_475; // @[util.scala 80:21]
  wire [31:0] _GEN_508 = wvalid ? _GEN_28 : _GEN_476; // @[util.scala 80:21]
  wire [31:0] _GEN_509 = wvalid ? _GEN_29 : _GEN_477; // @[util.scala 80:21]
  wire [31:0] _GEN_510 = wvalid ? _GEN_30 : _GEN_478; // @[util.scala 80:21]
  wire [31:0] _GEN_511 = wvalid ? _GEN_31 : _GEN_479; // @[util.scala 80:21]
  wire [31:0] _GEN_512 = wvalid ? _GEN_32 : _GEN_480; // @[util.scala 80:21]
  wire [31:0] _GEN_513 = wvalid ? _GEN_33 : _GEN_481; // @[util.scala 80:21]
  wire [31:0] _GEN_514 = wvalid ? _GEN_34 : _GEN_482; // @[util.scala 80:21]
  wire [31:0] _GEN_515 = wvalid ? _GEN_35 : _GEN_483; // @[util.scala 80:21]
  wire [31:0] _GEN_516 = wvalid ? _GEN_36 : _GEN_484; // @[util.scala 80:21]
  wire [31:0] _GEN_517 = wvalid ? _GEN_37 : _GEN_485; // @[util.scala 80:21]
  wire [31:0] _GEN_518 = wvalid ? _GEN_38 : _GEN_486; // @[util.scala 80:21]
  wire [31:0] _GEN_519 = wvalid ? _GEN_39 : _GEN_487; // @[util.scala 80:21]
  wire [31:0] _GEN_520 = wvalid ? _GEN_40 : _GEN_488; // @[util.scala 80:21]
  wire [31:0] _GEN_521 = wvalid ? _GEN_41 : _GEN_489; // @[util.scala 80:21]
  wire [31:0] _GEN_522 = wvalid ? _GEN_42 : _GEN_490; // @[util.scala 80:21]
  wire [31:0] _GEN_523 = wvalid ? _GEN_43 : _GEN_491; // @[util.scala 80:21]
  reg [4:0] eraddr; // @[util.scala 92:19]
  wire [31:0] _GEN_622 = 5'h1 == eraddr ? table_1 : table_0; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_623 = 5'h2 == eraddr ? table_2 : _GEN_622; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_624 = 5'h3 == eraddr ? table_3 : _GEN_623; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_625 = 5'h4 == eraddr ? table_4 : _GEN_624; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_626 = 5'h5 == eraddr ? table_5 : _GEN_625; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_627 = 5'h6 == eraddr ? table_6 : _GEN_626; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_628 = 5'h7 == eraddr ? table_7 : _GEN_627; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_629 = 5'h8 == eraddr ? table_8 : _GEN_628; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_630 = 5'h9 == eraddr ? table_9 : _GEN_629; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_631 = 5'ha == eraddr ? table_10 : _GEN_630; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_632 = 5'hb == eraddr ? table_11 : _GEN_631; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_633 = 5'hc == eraddr ? table_12 : _GEN_632; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_634 = 5'hd == eraddr ? table_13 : _GEN_633; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_635 = 5'he == eraddr ? table_14 : _GEN_634; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_636 = 5'hf == eraddr ? table_15 : _GEN_635; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_637 = 5'h10 == eraddr ? table_16 : _GEN_636; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_638 = 5'h11 == eraddr ? table_17 : _GEN_637; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_639 = 5'h12 == eraddr ? table_18 : _GEN_638; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_640 = 5'h13 == eraddr ? table_19 : _GEN_639; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_641 = 5'h14 == eraddr ? table_20 : _GEN_640; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_642 = 5'h15 == eraddr ? table_21 : _GEN_641; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_643 = 5'h16 == eraddr ? table_22 : _GEN_642; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_644 = 5'h17 == eraddr ? table_23 : _GEN_643; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_645 = 5'h18 == eraddr ? table_24 : _GEN_644; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_646 = 5'h19 == eraddr ? table_25 : _GEN_645; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_647 = 5'h1a == eraddr ? table_26 : _GEN_646; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_648 = 5'h1b == eraddr ? table_27 : _GEN_647; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_649 = 5'h1c == eraddr ? table_28 : _GEN_648; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_650 = 5'h1d == eraddr ? table_29 : _GEN_649; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_651 = 5'h1e == eraddr ? table_30 : _GEN_650; // @[util.scala 99:16 util.scala 99:16]
  assign io_data_0 = table_0; // @[util.scala 53:11]
  assign io_data_1 = table_1; // @[util.scala 53:11]
  assign io_data_2 = table_2; // @[util.scala 53:11]
  assign io_data_3 = table_3; // @[util.scala 53:11]
  assign io_data_4 = table_4; // @[util.scala 53:11]
  assign io_data_5 = table_5; // @[util.scala 53:11]
  assign io_data_6 = table_6; // @[util.scala 53:11]
  assign io_data_7 = table_7; // @[util.scala 53:11]
  assign io_data_8 = table_8; // @[util.scala 53:11]
  assign io_data_9 = table_9; // @[util.scala 53:11]
  assign io_data_10 = table_10; // @[util.scala 53:11]
  assign io_data_11 = table_11; // @[util.scala 53:11]
  assign io_data_12 = table_12; // @[util.scala 53:11]
  assign io_data_13 = table_13; // @[util.scala 53:11]
  assign config_awready = status == 3'h0; // @[util.scala 55:28]
  assign config_arready = status == 3'h0; // @[util.scala 56:28]
  assign config_wready = status == 3'h1; // @[util.scala 54:27]
  assign config_rdata = 5'h1f == eraddr ? table_31 : _GEN_651; // @[util.scala 99:16 util.scala 99:16]
  assign config_rvalid = status == 3'h5; // @[util.scala 57:27]
  assign config_bvalid = status == 3'h3; // @[util.scala 58:27]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 16:22]
      table_0 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h0 == io_wptr_1) begin // @[util.scala 73:23]
        table_0 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_0 <= _GEN_44;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_0 <= _GEN_44;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_0 <= _GEN_204;
    end else begin
      table_0 <= _GEN_492;
    end
    if (reset) begin // @[util.scala 16:22]
      table_1 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1 == io_wptr_1) begin // @[util.scala 73:23]
        table_1 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_1 <= _GEN_45;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_1 <= _GEN_45;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_1 <= _GEN_205;
    end else begin
      table_1 <= _GEN_493;
    end
    if (reset) begin // @[util.scala 16:22]
      table_2 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h2 == io_wptr_1) begin // @[util.scala 73:23]
        table_2 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_2 <= _GEN_46;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_2 <= _GEN_46;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_2 <= _GEN_206;
    end else begin
      table_2 <= _GEN_494;
    end
    if (reset) begin // @[util.scala 16:22]
      table_3 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h3 == io_wptr_1) begin // @[util.scala 73:23]
        table_3 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_3 <= _GEN_47;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_3 <= _GEN_47;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_3 <= _GEN_207;
    end else begin
      table_3 <= _GEN_495;
    end
    if (reset) begin // @[util.scala 16:22]
      table_4 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h4 == io_wptr_1) begin // @[util.scala 73:23]
        table_4 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_4 <= _GEN_48;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_4 <= _GEN_48;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_4 <= _GEN_208;
    end else begin
      table_4 <= _GEN_496;
    end
    if (reset) begin // @[util.scala 16:22]
      table_5 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h5 == io_wptr_1) begin // @[util.scala 73:23]
        table_5 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_5 <= _GEN_49;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_5 <= _GEN_49;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_5 <= _GEN_209;
    end else begin
      table_5 <= _GEN_497;
    end
    if (reset) begin // @[util.scala 16:22]
      table_6 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h6 == io_wptr_1) begin // @[util.scala 73:23]
        table_6 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_6 <= _GEN_50;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_6 <= _GEN_50;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_6 <= _GEN_210;
    end else begin
      table_6 <= _GEN_498;
    end
    if (reset) begin // @[util.scala 16:22]
      table_7 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h7 == io_wptr_1) begin // @[util.scala 73:23]
        table_7 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_7 <= _GEN_51;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_7 <= _GEN_51;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_7 <= _GEN_211;
    end else begin
      table_7 <= _GEN_499;
    end
    if (reset) begin // @[util.scala 16:22]
      table_8 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h8 == io_wptr_1) begin // @[util.scala 73:23]
        table_8 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_8 <= _GEN_52;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_8 <= _GEN_52;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_8 <= _GEN_212;
    end else begin
      table_8 <= _GEN_500;
    end
    if (reset) begin // @[util.scala 16:22]
      table_9 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h9 == io_wptr_1) begin // @[util.scala 73:23]
        table_9 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_9 <= _GEN_53;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_9 <= _GEN_53;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_9 <= _GEN_213;
    end else begin
      table_9 <= _GEN_501;
    end
    if (reset) begin // @[util.scala 16:22]
      table_10 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'ha == io_wptr_1) begin // @[util.scala 73:23]
        table_10 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_10 <= _GEN_54;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_10 <= _GEN_54;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_10 <= _GEN_214;
    end else begin
      table_10 <= _GEN_502;
    end
    if (reset) begin // @[util.scala 16:22]
      table_11 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hb == io_wptr_1) begin // @[util.scala 73:23]
        table_11 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_11 <= _GEN_55;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_11 <= _GEN_55;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_11 <= _GEN_215;
    end else begin
      table_11 <= _GEN_503;
    end
    if (reset) begin // @[util.scala 16:22]
      table_12 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hc == io_wptr_1) begin // @[util.scala 73:23]
        table_12 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_12 <= _GEN_56;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_12 <= _GEN_56;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_12 <= _GEN_216;
    end else begin
      table_12 <= _GEN_504;
    end
    if (reset) begin // @[util.scala 16:22]
      table_13 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hd == io_wptr_1) begin // @[util.scala 73:23]
        table_13 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_13 <= _GEN_57;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_13 <= _GEN_57;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_13 <= _GEN_217;
    end else begin
      table_13 <= _GEN_505;
    end
    if (reset) begin // @[util.scala 16:22]
      table_14 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'he == io_wptr_1) begin // @[util.scala 73:23]
        table_14 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_14 <= _GEN_58;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_14 <= _GEN_58;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_14 <= _GEN_218;
    end else begin
      table_14 <= _GEN_506;
    end
    if (reset) begin // @[util.scala 16:22]
      table_15 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hf == io_wptr_1) begin // @[util.scala 73:23]
        table_15 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_15 <= _GEN_59;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_15 <= _GEN_59;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_15 <= _GEN_219;
    end else begin
      table_15 <= _GEN_507;
    end
    if (reset) begin // @[util.scala 16:22]
      table_16 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h10 == io_wptr_1) begin // @[util.scala 73:23]
        table_16 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_16 <= _GEN_60;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_16 <= _GEN_60;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_16 <= _GEN_220;
    end else begin
      table_16 <= _GEN_508;
    end
    if (reset) begin // @[util.scala 16:22]
      table_17 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h11 == io_wptr_1) begin // @[util.scala 73:23]
        table_17 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_17 <= _GEN_61;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_17 <= _GEN_61;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_17 <= _GEN_221;
    end else begin
      table_17 <= _GEN_509;
    end
    if (reset) begin // @[util.scala 16:22]
      table_18 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h12 == io_wptr_1) begin // @[util.scala 73:23]
        table_18 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_18 <= _GEN_62;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_18 <= _GEN_62;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_18 <= _GEN_222;
    end else begin
      table_18 <= _GEN_510;
    end
    if (reset) begin // @[util.scala 16:22]
      table_19 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h13 == io_wptr_1) begin // @[util.scala 73:23]
        table_19 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_19 <= _GEN_63;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_19 <= _GEN_63;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_19 <= _GEN_223;
    end else begin
      table_19 <= _GEN_511;
    end
    if (reset) begin // @[util.scala 16:22]
      table_20 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h14 == io_wptr_1) begin // @[util.scala 73:23]
        table_20 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_20 <= _GEN_64;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_20 <= _GEN_64;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_20 <= _GEN_224;
    end else begin
      table_20 <= _GEN_512;
    end
    if (reset) begin // @[util.scala 16:22]
      table_21 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h15 == io_wptr_1) begin // @[util.scala 73:23]
        table_21 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_21 <= _GEN_65;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_21 <= _GEN_65;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_21 <= _GEN_225;
    end else begin
      table_21 <= _GEN_513;
    end
    if (reset) begin // @[util.scala 16:22]
      table_22 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h16 == io_wptr_1) begin // @[util.scala 73:23]
        table_22 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_22 <= _GEN_66;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_22 <= _GEN_66;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_22 <= _GEN_226;
    end else begin
      table_22 <= _GEN_514;
    end
    if (reset) begin // @[util.scala 16:22]
      table_23 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h17 == io_wptr_1) begin // @[util.scala 73:23]
        table_23 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_23 <= _GEN_67;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_23 <= _GEN_67;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_23 <= _GEN_227;
    end else begin
      table_23 <= _GEN_515;
    end
    if (reset) begin // @[util.scala 16:22]
      table_24 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h18 == io_wptr_1) begin // @[util.scala 73:23]
        table_24 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_24 <= _GEN_68;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_24 <= _GEN_68;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_24 <= _GEN_228;
    end else begin
      table_24 <= _GEN_516;
    end
    if (reset) begin // @[util.scala 16:22]
      table_25 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h19 == io_wptr_1) begin // @[util.scala 73:23]
        table_25 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_25 <= _GEN_69;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_25 <= _GEN_69;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_25 <= _GEN_229;
    end else begin
      table_25 <= _GEN_517;
    end
    if (reset) begin // @[util.scala 16:22]
      table_26 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1a == io_wptr_1) begin // @[util.scala 73:23]
        table_26 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_26 <= _GEN_70;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_26 <= _GEN_70;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_26 <= _GEN_230;
    end else begin
      table_26 <= _GEN_518;
    end
    if (reset) begin // @[util.scala 16:22]
      table_27 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1b == io_wptr_1) begin // @[util.scala 73:23]
        table_27 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_27 <= _GEN_71;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_27 <= _GEN_71;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_27 <= _GEN_231;
    end else begin
      table_27 <= _GEN_519;
    end
    if (reset) begin // @[util.scala 16:22]
      table_28 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1c == io_wptr_1) begin // @[util.scala 73:23]
        table_28 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_28 <= _GEN_72;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_28 <= _GEN_72;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_28 <= _GEN_232;
    end else begin
      table_28 <= _GEN_520;
    end
    if (reset) begin // @[util.scala 16:22]
      table_29 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1d == io_wptr_1) begin // @[util.scala 73:23]
        table_29 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_29 <= _GEN_73;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_29 <= _GEN_73;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_29 <= _GEN_233;
    end else begin
      table_29 <= _GEN_521;
    end
    if (reset) begin // @[util.scala 16:22]
      table_30 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1e == io_wptr_1) begin // @[util.scala 73:23]
        table_30 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_30 <= _GEN_74;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_30 <= _GEN_74;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_30 <= _GEN_234;
    end else begin
      table_30 <= _GEN_522;
    end
    if (reset) begin // @[util.scala 16:22]
      table_31 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1f == io_wptr_1) begin // @[util.scala 73:23]
        table_31 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_31 <= _GEN_75;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_31 <= _GEN_75;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_31 <= _GEN_235;
    end else begin
      table_31 <= _GEN_523;
    end
    if (reset) begin // @[util.scala 26:23]
      status <= 3'h0; // @[util.scala 26:23]
    end else if (status == 3'h0) begin // @[util.scala 28:28]
      if (config_awvalid) begin // @[util.scala 29:25]
        status <= 3'h1; // @[util.scala 30:14]
      end else if (config_arvalid) begin // @[util.scala 31:31]
        status <= 3'h4; // @[util.scala 32:14]
      end
    end else if (status == 3'h1) begin // @[util.scala 34:35]
      if (config_wvalid) begin // @[util.scala 35:24]
        status <= 3'h2; // @[util.scala 36:14]
      end
    end else if (status == 3'h2) begin // @[util.scala 38:34]
      status <= 3'h3; // @[util.scala 39:12]
    end else begin
      status <= _GEN_7;
    end
    if (config_awvalid & config_awready) begin // @[util.scala 66:41]
      ewaddr <= config_awaddr[6:2]; // @[util.scala 67:12]
    end
    if (config_arvalid & config_arready) begin // @[util.scala 93:41]
      eraddr <= config_araddr[6:2]; // @[util.scala 94:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  table_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  table_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  table_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  table_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  table_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  table_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  table_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  table_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  table_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  table_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  table_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  table_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  table_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  table_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  table_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  table_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  table_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  table_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  table_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  table_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  table_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  table_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  table_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  table_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  table_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  table_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  table_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  table_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  table_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  table_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  table_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  table_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  status = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  ewaddr = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  eraddr = _RAND_34[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module controller(
  input         clock,
  input         reset,
  output [31:0] io_data_0,
  output [31:0] io_data_1,
  output [31:0] io_data_2,
  output [31:0] io_data_3,
  output [31:0] io_data_4,
  output [31:0] io_data_5,
  output [31:0] io_data_6,
  output [31:0] io_data_7,
  output [31:0] io_data_8,
  output [31:0] io_data_9,
  output [31:0] io_data_10,
  output [31:0] io_data_11,
  input         io_fin_0,
  input         io_fin_1,
  input         io_fin_2,
  input         io_fin_3,
  input         io_fin_4,
  input         io_fin_5,
  input         io_fin_6,
  input         io_fin_7,
  input         io_fin_8,
  input         io_fin_9,
  input         io_fin_10,
  input         io_fin_11,
  input         io_fin_12,
  input         io_fin_13,
  input         io_fin_14,
  input         io_fin_15,
  output        io_signal,
  output        io_start,
  output [31:0] io_level,
  input  [31:0] io_unvisited_size,
  input  [63:0] io_traveled_edges,
  input  [63:0] io_config_awaddr,
  input         io_config_awvalid,
  output        io_config_awready,
  input  [63:0] io_config_araddr,
  input         io_config_arvalid,
  output        io_config_arready,
  input  [31:0] io_config_wdata,
  input         io_config_wvalid,
  output        io_config_wready,
  output [31:0] io_config_rdata,
  output        io_config_rvalid,
  input         io_config_rready,
  output        io_config_bvalid,
  input         io_config_bready,
  output        io_flush_cache,
  input         io_flush_cache_end,
  input         io_signal_ack
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire  controls_clock; // @[BFS.scala 1430:24]
  wire  controls_reset; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_0; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_1; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_2; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_3; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_4; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_5; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_6; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_7; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_8; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_9; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_10; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_11; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_12; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_data_13; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_dataIn_0; // @[BFS.scala 1430:24]
  wire [31:0] controls_io_dataIn_1; // @[BFS.scala 1430:24]
  wire  controls_io_writeFlag_0; // @[BFS.scala 1430:24]
  wire  controls_io_writeFlag_1; // @[BFS.scala 1430:24]
  wire [4:0] controls_io_wptr_0; // @[BFS.scala 1430:24]
  wire [4:0] controls_io_wptr_1; // @[BFS.scala 1430:24]
  wire [63:0] controls_config_awaddr; // @[BFS.scala 1430:24]
  wire  controls_config_awvalid; // @[BFS.scala 1430:24]
  wire  controls_config_awready; // @[BFS.scala 1430:24]
  wire [63:0] controls_config_araddr; // @[BFS.scala 1430:24]
  wire  controls_config_arvalid; // @[BFS.scala 1430:24]
  wire  controls_config_arready; // @[BFS.scala 1430:24]
  wire [31:0] controls_config_wdata; // @[BFS.scala 1430:24]
  wire  controls_config_wvalid; // @[BFS.scala 1430:24]
  wire  controls_config_wready; // @[BFS.scala 1430:24]
  wire [31:0] controls_config_rdata; // @[BFS.scala 1430:24]
  wire  controls_config_rvalid; // @[BFS.scala 1430:24]
  wire  controls_config_rready; // @[BFS.scala 1430:24]
  wire  controls_config_bvalid; // @[BFS.scala 1430:24]
  wire  controls_config_bready; // @[BFS.scala 1430:24]
    (*dont_touch = "true" *)reg [31:0] level; // @[BFS.scala 1431:22]
  reg [2:0] status; // @[BFS.scala 1441:23]
  wire  start = controls_io_data_0[0] & ~controls_io_data_0[1]; // @[BFS.scala 1442:38]
  reg  FIN_0; // @[BFS.scala 1443:20]
  reg  FIN_1; // @[BFS.scala 1443:20]
  reg  FIN_2; // @[BFS.scala 1443:20]
  reg  FIN_3; // @[BFS.scala 1443:20]
  reg  FIN_4; // @[BFS.scala 1443:20]
  reg  FIN_5; // @[BFS.scala 1443:20]
  reg  FIN_6; // @[BFS.scala 1443:20]
  reg  FIN_7; // @[BFS.scala 1443:20]
  reg  FIN_8; // @[BFS.scala 1443:20]
  reg  FIN_9; // @[BFS.scala 1443:20]
  reg  FIN_10; // @[BFS.scala 1443:20]
  reg  FIN_11; // @[BFS.scala 1443:20]
  reg  FIN_12; // @[BFS.scala 1443:20]
  reg  FIN_13; // @[BFS.scala 1443:20]
  reg  FIN_14; // @[BFS.scala 1443:20]
  reg  FIN_15; // @[BFS.scala 1443:20]
  wire [63:0] _new_tep_T = {controls_io_data_12,controls_io_data_13}; // @[Cat.scala 30:58]
  wire [63:0] new_tep = _new_tep_T + io_traveled_edges; // @[BFS.scala 1444:65]
  reg [63:0] counterValue; // @[BFS.scala 1445:29]
  wire  _controls_io_writeFlag_0_T = status == 3'h3; // @[BFS.scala 1448:38]
  wire  _controls_io_writeFlag_0_T_1 = status == 3'h2; // @[BFS.scala 1448:59]
  wire  _controls_io_writeFlag_0_T_3 = status == 3'h2 & io_signal_ack; // @[BFS.scala 1448:70]
  wire  _controls_io_writeFlag_0_T_5 = status == 3'h6; // @[BFS.scala 1448:108]
  wire [3:0] _controls_io_wptr_0_T_3 = _controls_io_writeFlag_0_T_1 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_0_T_4 = _controls_io_writeFlag_0_T_5 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_0_T_6 = _controls_io_wptr_0_T_3 | _controls_io_wptr_0_T_4; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_5 = _controls_io_writeFlag_0_T_1 ? new_tep[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_6 = _controls_io_writeFlag_0_T_5 ? counterValue[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [1:0] _controls_io_dataIn_0_T_7 = _controls_io_writeFlag_0_T ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_8 = _controls_io_dataIn_0_T_5 | _controls_io_dataIn_0_T_6; // @[Mux.scala 27:72]
  wire [31:0] _GEN_44 = {{30'd0}, _controls_io_dataIn_0_T_7}; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_1_T_1 = _controls_io_writeFlag_0_T_1 ? 4'hd : 4'hf; // @[BFS.scala 1460:29]
  wire [31:0] _controls_io_dataIn_1_T_4 = _controls_io_writeFlag_0_T_1 ? new_tep[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_1_T_5 = _controls_io_writeFlag_0_T_5 ? counterValue[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1 = status == 3'h0 & start; // @[BFS.scala 1466:28]
  wire  _T_2 = status == 3'h4; // @[BFS.scala 1468:21]
  wire [2:0] _GEN_0 = io_unvisited_size == 32'h0 ? 3'h6 : 3'h1; // @[BFS.scala 1473:36 BFS.scala 1474:14 BFS.scala 1476:14]
  wire [2:0] _GEN_1 = _controls_io_writeFlag_0_T_5 ? 3'h5 : status; // @[BFS.scala 1480:40 BFS.scala 1481:12 BFS.scala 1441:23]
  wire [2:0] _GEN_2 = status == 3'h5 & io_flush_cache_end ? 3'h3 : _GEN_1; // @[BFS.scala 1478:62 BFS.scala 1479:12]
  wire [2:0] _GEN_3 = _controls_io_writeFlag_0_T_3 ? _GEN_0 : _GEN_2; // @[BFS.scala 1472:60]
  wire  _GEN_7 = io_fin_0 | FIN_0; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_9 = io_fin_1 | FIN_1; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_11 = io_fin_2 | FIN_2; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_13 = io_fin_3 | FIN_3; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_15 = io_fin_4 | FIN_4; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_17 = io_fin_5 | FIN_5; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_19 = io_fin_6 | FIN_6; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_21 = io_fin_7 | FIN_7; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_23 = io_fin_8 | FIN_8; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_25 = io_fin_9 | FIN_9; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_27 = io_fin_10 | FIN_10; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_29 = io_fin_11 | FIN_11; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_31 = io_fin_12 | FIN_12; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_33 = io_fin_13 | FIN_13; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_35 = io_fin_14 | FIN_14; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire  _GEN_37 = io_fin_15 | FIN_15; // @[BFS.scala 1490:28 BFS.scala 1491:11 BFS.scala 1443:20]
  wire [31:0] _level_T_1 = level + 32'h1; // @[BFS.scala 1497:20]
  wire  global_start = _controls_io_writeFlag_0_T_3 & level == 32'hffffffff; // @[BFS.scala 1502:68]
  wire [63:0] _counterValue_T_1 = counterValue + 64'h1; // @[BFS.scala 1506:34]
  reg [63:0] performanceValue_0; // @[BFS.scala 1509:33]
  LookupTable controls ( // @[BFS.scala 1430:24]
    .clock(controls_clock),
    .reset(controls_reset),
    .io_data_0(controls_io_data_0),
    .io_data_1(controls_io_data_1),
    .io_data_2(controls_io_data_2),
    .io_data_3(controls_io_data_3),
    .io_data_4(controls_io_data_4),
    .io_data_5(controls_io_data_5),
    .io_data_6(controls_io_data_6),
    .io_data_7(controls_io_data_7),
    .io_data_8(controls_io_data_8),
    .io_data_9(controls_io_data_9),
    .io_data_10(controls_io_data_10),
    .io_data_11(controls_io_data_11),
    .io_data_12(controls_io_data_12),
    .io_data_13(controls_io_data_13),
    .io_dataIn_0(controls_io_dataIn_0),
    .io_dataIn_1(controls_io_dataIn_1),
    .io_writeFlag_0(controls_io_writeFlag_0),
    .io_writeFlag_1(controls_io_writeFlag_1),
    .io_wptr_0(controls_io_wptr_0),
    .io_wptr_1(controls_io_wptr_1),
    .config_awaddr(controls_config_awaddr),
    .config_awvalid(controls_config_awvalid),
    .config_awready(controls_config_awready),
    .config_araddr(controls_config_araddr),
    .config_arvalid(controls_config_arvalid),
    .config_arready(controls_config_arready),
    .config_wdata(controls_config_wdata),
    .config_wvalid(controls_config_wvalid),
    .config_wready(controls_config_wready),
    .config_rdata(controls_config_rdata),
    .config_rvalid(controls_config_rvalid),
    .config_rready(controls_config_rready),
    .config_bvalid(controls_config_bvalid),
    .config_bready(controls_config_bready)
  );
  assign io_data_0 = controls_io_data_0; // @[BFS.scala 1522:11]
  assign io_data_1 = controls_io_data_1; // @[BFS.scala 1522:11]
  assign io_data_2 = controls_io_data_2; // @[BFS.scala 1522:11]
  assign io_data_3 = controls_io_data_3; // @[BFS.scala 1522:11]
  assign io_data_4 = controls_io_data_4; // @[BFS.scala 1522:11]
  assign io_data_5 = controls_io_data_5; // @[BFS.scala 1522:11]
  assign io_data_6 = controls_io_data_6; // @[BFS.scala 1522:11]
  assign io_data_7 = controls_io_data_7; // @[BFS.scala 1522:11]
  assign io_data_8 = controls_io_data_8; // @[BFS.scala 1522:11]
  assign io_data_9 = controls_io_data_9; // @[BFS.scala 1522:11]
  assign io_data_10 = controls_io_data_10; // @[BFS.scala 1522:11]
  assign io_data_11 = controls_io_data_11; // @[BFS.scala 1522:11]
  assign io_signal = _T_2 | _controls_io_writeFlag_0_T_1 & io_unvisited_size != 32'h0; // @[BFS.scala 1521:36]
  assign io_start = status == 3'h4; // @[BFS.scala 1524:22]
  assign io_level = level; // @[BFS.scala 1523:12]
  assign io_config_awready = controls_config_awready; // @[BFS.scala 1447:19]
  assign io_config_arready = controls_config_arready; // @[BFS.scala 1447:19]
  assign io_config_wready = controls_config_wready; // @[BFS.scala 1447:19]
  assign io_config_rdata = controls_config_rdata; // @[BFS.scala 1447:19]
  assign io_config_rvalid = controls_config_rvalid; // @[BFS.scala 1447:19]
  assign io_config_bvalid = controls_config_bvalid; // @[BFS.scala 1447:19]
  assign io_flush_cache = status == 3'h5; // @[BFS.scala 1525:28]
  assign controls_clock = clock;
  assign controls_reset = reset;
  assign controls_io_dataIn_0 = _controls_io_dataIn_0_T_8 | _GEN_44; // @[Mux.scala 27:72]
  assign controls_io_dataIn_1 = _controls_io_dataIn_1_T_4 | _controls_io_dataIn_1_T_5; // @[Mux.scala 27:72]
  assign controls_io_writeFlag_0 = status == 3'h3 | status == 3'h2 & io_signal_ack | status == 3'h6; // @[BFS.scala 1448:99]
  assign controls_io_writeFlag_1 = _controls_io_writeFlag_0_T_3 | _controls_io_writeFlag_0_T_5; // @[BFS.scala 1459:79]
  assign controls_io_wptr_0 = {{1'd0}, _controls_io_wptr_0_T_6}; // @[Mux.scala 27:72]
  assign controls_io_wptr_1 = {{1'd0}, _controls_io_wptr_1_T_1}; // @[BFS.scala 1460:29]
  assign controls_config_awaddr = io_config_awaddr; // @[BFS.scala 1447:19]
  assign controls_config_awvalid = io_config_awvalid; // @[BFS.scala 1447:19]
  assign controls_config_araddr = io_config_araddr; // @[BFS.scala 1447:19]
  assign controls_config_arvalid = io_config_arvalid; // @[BFS.scala 1447:19]
  assign controls_config_wdata = io_config_wdata; // @[BFS.scala 1447:19]
  assign controls_config_wvalid = io_config_wvalid; // @[BFS.scala 1447:19]
  assign controls_config_rready = io_config_rready; // @[BFS.scala 1447:19]
  assign controls_config_bready = io_config_bready; // @[BFS.scala 1447:19]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1431:22]
      level <= 32'h0; // @[BFS.scala 1431:22]
    end else if (_controls_io_writeFlag_0_T_3) begin // @[BFS.scala 1496:54]
      level <= _level_T_1; // @[BFS.scala 1497:11]
    end else if (_T_1) begin // @[BFS.scala 1498:43]
      level <= 32'hffffffff; // @[BFS.scala 1499:11]
    end
    if (reset) begin // @[BFS.scala 1441:23]
      status <= 3'h0; // @[BFS.scala 1441:23]
    end else if (status == 3'h0 & start) begin // @[BFS.scala 1466:37]
      status <= 3'h4; // @[BFS.scala 1467:12]
    end else if (status == 3'h4) begin // @[BFS.scala 1468:34]
      status <= 3'h1; // @[BFS.scala 1469:12]
    end else if (status == 3'h1 & (FIN_0 & FIN_1 & FIN_2 & FIN_3 & FIN_4 & FIN_5 & FIN_6 & FIN_7 & FIN_8 & FIN_9 &
      FIN_10 & FIN_11 & FIN_12 & FIN_13 & FIN_14 & FIN_15)) begin // @[BFS.scala 1470:51]
      status <= 3'h2; // @[BFS.scala 1471:12]
    end else begin
      status <= _GEN_3;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_0 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_0 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_0 <= _GEN_7;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_1 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_1 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_1 <= _GEN_9;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_2 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_2 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_2 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_3 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_3 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_3 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_4 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_4 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_4 <= _GEN_15;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_5 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_5 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_5 <= _GEN_17;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_6 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_6 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_6 <= _GEN_19;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_7 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_7 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_7 <= _GEN_21;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_8 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_8 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_8 <= _GEN_23;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_9 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_9 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_9 <= _GEN_25;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_10 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_10 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_10 <= _GEN_27;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_11 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_11 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_11 <= _GEN_29;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_12 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_12 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_12 <= _GEN_31;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_13 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_13 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_13 <= _GEN_33;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_14 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_14 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_14 <= _GEN_35;
    end
    if (reset) begin // @[BFS.scala 1443:20]
      FIN_15 <= 1'h0; // @[BFS.scala 1443:20]
    end else if (io_signal) begin // @[BFS.scala 1488:22]
      FIN_15 <= 1'h0; // @[BFS.scala 1489:11]
    end else begin
      FIN_15 <= _GEN_37;
    end
    if (reset) begin // @[BFS.scala 1445:29]
      counterValue <= 64'h0; // @[BFS.scala 1445:29]
    end else if (global_start) begin // @[BFS.scala 1503:22]
      counterValue <= 64'h0; // @[BFS.scala 1504:18]
    end else begin
      counterValue <= _counterValue_T_1; // @[BFS.scala 1506:18]
    end
    if (reset) begin // @[BFS.scala 1509:33]
      performanceValue_0 <= 64'h0; // @[BFS.scala 1509:33]
    end else if (global_start) begin // @[BFS.scala 1513:26]
      performanceValue_0 <= 64'h0; // @[BFS.scala 1514:29]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  level = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  status = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  FIN_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIN_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  FIN_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  FIN_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  FIN_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  FIN_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  FIN_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  FIN_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  FIN_8 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  FIN_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  FIN_10 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  FIN_11 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  FIN_12 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  FIN_13 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  FIN_14 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  FIN_15 = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  counterValue = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  performanceValue_0 = _RAND_19[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multi_channel_fifo(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [31:0]  io_in_bits_0_tdata,
  input          io_in_bits_0_tkeep,
  input  [31:0]  io_in_bits_1_tdata,
  input          io_in_bits_1_tkeep,
  input  [31:0]  io_in_bits_2_tdata,
  input          io_in_bits_2_tkeep,
  input  [31:0]  io_in_bits_3_tdata,
  input          io_in_bits_3_tkeep,
  input  [31:0]  io_in_bits_4_tdata,
  input          io_in_bits_4_tkeep,
  input  [31:0]  io_in_bits_5_tdata,
  input          io_in_bits_5_tkeep,
  input  [31:0]  io_in_bits_6_tdata,
  input          io_in_bits_6_tkeep,
  input  [31:0]  io_in_bits_7_tdata,
  input          io_in_bits_7_tkeep,
  input  [31:0]  io_in_bits_8_tdata,
  input          io_in_bits_8_tkeep,
  input  [31:0]  io_in_bits_9_tdata,
  input          io_in_bits_9_tkeep,
  input  [31:0]  io_in_bits_10_tdata,
  input          io_in_bits_10_tkeep,
  input  [31:0]  io_in_bits_11_tdata,
  input          io_in_bits_11_tkeep,
  input  [31:0]  io_in_bits_12_tdata,
  input          io_in_bits_12_tkeep,
  input  [31:0]  io_in_bits_13_tdata,
  input          io_in_bits_13_tkeep,
  input  [31:0]  io_in_bits_14_tdata,
  input          io_in_bits_14_tkeep,
  input  [31:0]  io_in_bits_15_tdata,
  input          io_in_bits_15_tkeep,
  output         io_out_almost_full,
  input  [511:0] io_out_din,
  input          io_out_wr_en,
  output [511:0] io_out_dout,
  input          io_out_rd_en,
  output [13:0]  io_out_data_count,
  output         io_out_valid,
  input          io_is_current_tier
);
  wire  collector_fifos_0_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_0_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_0_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_0_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_0_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_0_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_0_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_0_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_0_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_0_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_1_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_1_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_1_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_1_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_1_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_1_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_1_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_1_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_1_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_1_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_2_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_2_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_2_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_2_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_2_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_2_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_2_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_2_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_2_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_2_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_3_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_3_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_3_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_3_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_3_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_3_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_3_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_3_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_3_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_3_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_4_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_4_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_4_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_4_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_4_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_4_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_4_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_4_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_4_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_4_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_5_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_5_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_5_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_5_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_5_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_5_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_5_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_5_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_5_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_5_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_6_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_6_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_6_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_6_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_6_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_6_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_6_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_6_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_6_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_6_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_7_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_7_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_7_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_7_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_7_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_7_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_7_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_7_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_7_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_7_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_8_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_8_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_8_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_8_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_8_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_8_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_8_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_8_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_8_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_8_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_9_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_9_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_9_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_9_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_9_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_9_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_9_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_9_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_9_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_9_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_10_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_10_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_10_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_10_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_10_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_10_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_10_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_10_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_10_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_10_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_11_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_11_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_11_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_11_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_11_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_11_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_11_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_11_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_11_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_11_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_12_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_12_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_12_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_12_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_12_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_12_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_12_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_12_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_12_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_12_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_13_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_13_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_13_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_13_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_13_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_13_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_13_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_13_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_13_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_13_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_14_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_14_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_14_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_14_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_14_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_14_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_14_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_14_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_14_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_14_valid; // @[BFS.scala 1134:16]
  wire  collector_fifos_15_full; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_15_din; // @[BFS.scala 1134:16]
  wire  collector_fifos_15_wr_en; // @[BFS.scala 1134:16]
  wire  collector_fifos_15_empty; // @[BFS.scala 1134:16]
  wire [31:0] collector_fifos_15_dout; // @[BFS.scala 1134:16]
  wire  collector_fifos_15_rd_en; // @[BFS.scala 1134:16]
  wire [9:0] collector_fifos_15_data_count; // @[BFS.scala 1134:16]
  wire  collector_fifos_15_clk; // @[BFS.scala 1134:16]
  wire  collector_fifos_15_srst; // @[BFS.scala 1134:16]
  wire  collector_fifos_15_valid; // @[BFS.scala 1134:16]
  wire  _io_in_ready_T_15 = ~collector_fifos_15_full; // @[BFS.scala 1137:67]
  wire [31:0] collector_data_1 = collector_fifos_1_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_0 = collector_fifos_0_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_3 = collector_fifos_3_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_2 = collector_fifos_2_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_5 = collector_fifos_5_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_4 = collector_fifos_4_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_7 = collector_fifos_7_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_6 = collector_fifos_6_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [255:0] io_out_dout_lo = {collector_data_7,collector_data_6,collector_data_5,collector_data_4,collector_data_3,
    collector_data_2,collector_data_1,collector_data_0}; // @[BFS.scala 1150:39]
  wire [31:0] collector_data_9 = collector_fifos_9_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_8 = collector_fifos_8_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_11 = collector_fifos_11_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_10 = collector_fifos_10_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_13 = collector_fifos_13_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_12 = collector_fifos_12_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_15 = collector_fifos_15_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [31:0] collector_data_14 = collector_fifos_14_dout; // @[BFS.scala 1136:28 BFS.scala 1142:25]
  wire [255:0] io_out_dout_hi = {collector_data_15,collector_data_14,collector_data_13,collector_data_12,
    collector_data_11,collector_data_10,collector_data_9,collector_data_8}; // @[BFS.scala 1150:39]
  wire [13:0] _io_out_data_count_WIRE = {{4'd0}, collector_fifos_0_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_WIRE_1 = {{4'd0}, collector_fifos_1_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_1 = _io_out_data_count_WIRE + _io_out_data_count_WIRE_1; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_2 = {{4'd0}, collector_fifos_2_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_3 = _io_out_data_count_T_1 + _io_out_data_count_WIRE_2; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_3 = {{4'd0}, collector_fifos_3_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_5 = _io_out_data_count_T_3 + _io_out_data_count_WIRE_3; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_4 = {{4'd0}, collector_fifos_4_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_7 = _io_out_data_count_T_5 + _io_out_data_count_WIRE_4; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_5 = {{4'd0}, collector_fifos_5_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_9 = _io_out_data_count_T_7 + _io_out_data_count_WIRE_5; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_6 = {{4'd0}, collector_fifos_6_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_11 = _io_out_data_count_T_9 + _io_out_data_count_WIRE_6; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_7 = {{4'd0}, collector_fifos_7_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_13 = _io_out_data_count_T_11 + _io_out_data_count_WIRE_7; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_8 = {{4'd0}, collector_fifos_8_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_15 = _io_out_data_count_T_13 + _io_out_data_count_WIRE_8; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_9 = {{4'd0}, collector_fifos_9_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_17 = _io_out_data_count_T_15 + _io_out_data_count_WIRE_9; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_10 = {{4'd0}, collector_fifos_10_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_19 = _io_out_data_count_T_17 + _io_out_data_count_WIRE_10; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_11 = {{4'd0}, collector_fifos_11_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_21 = _io_out_data_count_T_19 + _io_out_data_count_WIRE_11; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_12 = {{4'd0}, collector_fifos_12_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_23 = _io_out_data_count_T_21 + _io_out_data_count_WIRE_12; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_13 = {{4'd0}, collector_fifos_13_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_25 = _io_out_data_count_T_23 + _io_out_data_count_WIRE_13; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_14 = {{4'd0}, collector_fifos_14_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire [13:0] _io_out_data_count_T_27 = _io_out_data_count_T_25 + _io_out_data_count_WIRE_14; // @[BFS.scala 1153:13]
  wire [13:0] _io_out_data_count_WIRE_15 = {{4'd0}, collector_fifos_15_data_count}; // @[BFS.scala 1152:34 BFS.scala 1152:34]
  wire  _io_out_almost_full_T = collector_fifos_0_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_1 = collector_fifos_1_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_2 = collector_fifos_2_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_3 = collector_fifos_3_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_4 = collector_fifos_4_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_5 = collector_fifos_5_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_6 = collector_fifos_6_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_7 = collector_fifos_7_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_8 = collector_fifos_8_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_9 = collector_fifos_9_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_10 = collector_fifos_10_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_11 = collector_fifos_11_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_12 = collector_fifos_12_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_13 = collector_fifos_13_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_14 = collector_fifos_14_data_count > 10'h100; // @[BFS.scala 1155:27]
  wire  _io_out_almost_full_T_15 = collector_fifos_15_data_count > 10'h100; // @[BFS.scala 1155:27]
  collector_fifo_0 collector_fifos_0 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_0_full),
    .din(collector_fifos_0_din),
    .wr_en(collector_fifos_0_wr_en),
    .empty(collector_fifos_0_empty),
    .dout(collector_fifos_0_dout),
    .rd_en(collector_fifos_0_rd_en),
    .data_count(collector_fifos_0_data_count),
    .clk(collector_fifos_0_clk),
    .srst(collector_fifos_0_srst),
    .valid(collector_fifos_0_valid)
  );
  collector_fifo_0 collector_fifos_1 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_1_full),
    .din(collector_fifos_1_din),
    .wr_en(collector_fifos_1_wr_en),
    .empty(collector_fifos_1_empty),
    .dout(collector_fifos_1_dout),
    .rd_en(collector_fifos_1_rd_en),
    .data_count(collector_fifos_1_data_count),
    .clk(collector_fifos_1_clk),
    .srst(collector_fifos_1_srst),
    .valid(collector_fifos_1_valid)
  );
  collector_fifo_0 collector_fifos_2 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_2_full),
    .din(collector_fifos_2_din),
    .wr_en(collector_fifos_2_wr_en),
    .empty(collector_fifos_2_empty),
    .dout(collector_fifos_2_dout),
    .rd_en(collector_fifos_2_rd_en),
    .data_count(collector_fifos_2_data_count),
    .clk(collector_fifos_2_clk),
    .srst(collector_fifos_2_srst),
    .valid(collector_fifos_2_valid)
  );
  collector_fifo_0 collector_fifos_3 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_3_full),
    .din(collector_fifos_3_din),
    .wr_en(collector_fifos_3_wr_en),
    .empty(collector_fifos_3_empty),
    .dout(collector_fifos_3_dout),
    .rd_en(collector_fifos_3_rd_en),
    .data_count(collector_fifos_3_data_count),
    .clk(collector_fifos_3_clk),
    .srst(collector_fifos_3_srst),
    .valid(collector_fifos_3_valid)
  );
  collector_fifo_0 collector_fifos_4 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_4_full),
    .din(collector_fifos_4_din),
    .wr_en(collector_fifos_4_wr_en),
    .empty(collector_fifos_4_empty),
    .dout(collector_fifos_4_dout),
    .rd_en(collector_fifos_4_rd_en),
    .data_count(collector_fifos_4_data_count),
    .clk(collector_fifos_4_clk),
    .srst(collector_fifos_4_srst),
    .valid(collector_fifos_4_valid)
  );
  collector_fifo_0 collector_fifos_5 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_5_full),
    .din(collector_fifos_5_din),
    .wr_en(collector_fifos_5_wr_en),
    .empty(collector_fifos_5_empty),
    .dout(collector_fifos_5_dout),
    .rd_en(collector_fifos_5_rd_en),
    .data_count(collector_fifos_5_data_count),
    .clk(collector_fifos_5_clk),
    .srst(collector_fifos_5_srst),
    .valid(collector_fifos_5_valid)
  );
  collector_fifo_0 collector_fifos_6 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_6_full),
    .din(collector_fifos_6_din),
    .wr_en(collector_fifos_6_wr_en),
    .empty(collector_fifos_6_empty),
    .dout(collector_fifos_6_dout),
    .rd_en(collector_fifos_6_rd_en),
    .data_count(collector_fifos_6_data_count),
    .clk(collector_fifos_6_clk),
    .srst(collector_fifos_6_srst),
    .valid(collector_fifos_6_valid)
  );
  collector_fifo_0 collector_fifos_7 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_7_full),
    .din(collector_fifos_7_din),
    .wr_en(collector_fifos_7_wr_en),
    .empty(collector_fifos_7_empty),
    .dout(collector_fifos_7_dout),
    .rd_en(collector_fifos_7_rd_en),
    .data_count(collector_fifos_7_data_count),
    .clk(collector_fifos_7_clk),
    .srst(collector_fifos_7_srst),
    .valid(collector_fifos_7_valid)
  );
  collector_fifo_0 collector_fifos_8 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_8_full),
    .din(collector_fifos_8_din),
    .wr_en(collector_fifos_8_wr_en),
    .empty(collector_fifos_8_empty),
    .dout(collector_fifos_8_dout),
    .rd_en(collector_fifos_8_rd_en),
    .data_count(collector_fifos_8_data_count),
    .clk(collector_fifos_8_clk),
    .srst(collector_fifos_8_srst),
    .valid(collector_fifos_8_valid)
  );
  collector_fifo_0 collector_fifos_9 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_9_full),
    .din(collector_fifos_9_din),
    .wr_en(collector_fifos_9_wr_en),
    .empty(collector_fifos_9_empty),
    .dout(collector_fifos_9_dout),
    .rd_en(collector_fifos_9_rd_en),
    .data_count(collector_fifos_9_data_count),
    .clk(collector_fifos_9_clk),
    .srst(collector_fifos_9_srst),
    .valid(collector_fifos_9_valid)
  );
  collector_fifo_0 collector_fifos_10 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_10_full),
    .din(collector_fifos_10_din),
    .wr_en(collector_fifos_10_wr_en),
    .empty(collector_fifos_10_empty),
    .dout(collector_fifos_10_dout),
    .rd_en(collector_fifos_10_rd_en),
    .data_count(collector_fifos_10_data_count),
    .clk(collector_fifos_10_clk),
    .srst(collector_fifos_10_srst),
    .valid(collector_fifos_10_valid)
  );
  collector_fifo_0 collector_fifos_11 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_11_full),
    .din(collector_fifos_11_din),
    .wr_en(collector_fifos_11_wr_en),
    .empty(collector_fifos_11_empty),
    .dout(collector_fifos_11_dout),
    .rd_en(collector_fifos_11_rd_en),
    .data_count(collector_fifos_11_data_count),
    .clk(collector_fifos_11_clk),
    .srst(collector_fifos_11_srst),
    .valid(collector_fifos_11_valid)
  );
  collector_fifo_0 collector_fifos_12 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_12_full),
    .din(collector_fifos_12_din),
    .wr_en(collector_fifos_12_wr_en),
    .empty(collector_fifos_12_empty),
    .dout(collector_fifos_12_dout),
    .rd_en(collector_fifos_12_rd_en),
    .data_count(collector_fifos_12_data_count),
    .clk(collector_fifos_12_clk),
    .srst(collector_fifos_12_srst),
    .valid(collector_fifos_12_valid)
  );
  collector_fifo_0 collector_fifos_13 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_13_full),
    .din(collector_fifos_13_din),
    .wr_en(collector_fifos_13_wr_en),
    .empty(collector_fifos_13_empty),
    .dout(collector_fifos_13_dout),
    .rd_en(collector_fifos_13_rd_en),
    .data_count(collector_fifos_13_data_count),
    .clk(collector_fifos_13_clk),
    .srst(collector_fifos_13_srst),
    .valid(collector_fifos_13_valid)
  );
  collector_fifo_0 collector_fifos_14 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_14_full),
    .din(collector_fifos_14_din),
    .wr_en(collector_fifos_14_wr_en),
    .empty(collector_fifos_14_empty),
    .dout(collector_fifos_14_dout),
    .rd_en(collector_fifos_14_rd_en),
    .data_count(collector_fifos_14_data_count),
    .clk(collector_fifos_14_clk),
    .srst(collector_fifos_14_srst),
    .valid(collector_fifos_14_valid)
  );
  collector_fifo_0 collector_fifos_15 ( // @[BFS.scala 1134:16]
    .full(collector_fifos_15_full),
    .din(collector_fifos_15_din),
    .wr_en(collector_fifos_15_wr_en),
    .empty(collector_fifos_15_empty),
    .dout(collector_fifos_15_dout),
    .rd_en(collector_fifos_15_rd_en),
    .data_count(collector_fifos_15_data_count),
    .clk(collector_fifos_15_clk),
    .srst(collector_fifos_15_srst),
    .valid(collector_fifos_15_valid)
  );
  assign io_in_ready = ~collector_fifos_0_full & ~collector_fifos_1_full & ~collector_fifos_2_full & ~
    collector_fifos_3_full & ~collector_fifos_4_full & ~collector_fifos_5_full & ~collector_fifos_6_full & ~
    collector_fifos_7_full & ~collector_fifos_8_full & ~collector_fifos_9_full & ~collector_fifos_10_full & ~
    collector_fifos_11_full & ~collector_fifos_12_full & ~collector_fifos_13_full & ~collector_fifos_14_full &
    _io_in_ready_T_15; // @[BFS.scala 1137:88]
  assign io_out_almost_full = _io_out_almost_full_T & _io_out_almost_full_T_1 & _io_out_almost_full_T_2 &
    _io_out_almost_full_T_3 & _io_out_almost_full_T_4 & _io_out_almost_full_T_5 & _io_out_almost_full_T_6 &
    _io_out_almost_full_T_7 & _io_out_almost_full_T_8 & _io_out_almost_full_T_9 & _io_out_almost_full_T_10 &
    _io_out_almost_full_T_11 & _io_out_almost_full_T_12 & _io_out_almost_full_T_13 & _io_out_almost_full_T_14 &
    _io_out_almost_full_T_15; // @[BFS.scala 1156:13]
  assign io_out_dout = {io_out_dout_hi,io_out_dout_lo}; // @[BFS.scala 1150:39]
  assign io_out_data_count = _io_out_data_count_T_27 + _io_out_data_count_WIRE_15; // @[BFS.scala 1153:13]
  assign io_out_valid = collector_fifos_0_valid | collector_fifos_1_valid | collector_fifos_2_valid |
    collector_fifos_3_valid | collector_fifos_4_valid | collector_fifos_5_valid | collector_fifos_6_valid |
    collector_fifos_7_valid | collector_fifos_8_valid | collector_fifos_9_valid | collector_fifos_10_valid |
    collector_fifos_11_valid | collector_fifos_12_valid | collector_fifos_13_valid | collector_fifos_14_valid |
    collector_fifos_15_valid; // @[BFS.scala 1149:80]
  assign collector_fifos_0_din = io_is_current_tier ? io_out_din[31:0] : io_in_bits_0_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_0_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_0_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_0_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_0_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_0_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_1_din = io_is_current_tier ? io_out_din[63:32] : io_in_bits_1_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_1_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_1_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_1_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_1_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_1_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_2_din = io_is_current_tier ? io_out_din[95:64] : io_in_bits_2_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_2_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_2_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_2_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_2_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_2_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_3_din = io_is_current_tier ? io_out_din[127:96] : io_in_bits_3_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_3_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_3_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_3_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_3_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_3_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_4_din = io_is_current_tier ? io_out_din[159:128] : io_in_bits_4_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_4_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_4_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_4_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_4_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_4_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_5_din = io_is_current_tier ? io_out_din[191:160] : io_in_bits_5_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_5_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_5_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_5_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_5_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_5_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_6_din = io_is_current_tier ? io_out_din[223:192] : io_in_bits_6_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_6_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_6_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_6_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_6_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_6_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_7_din = io_is_current_tier ? io_out_din[255:224] : io_in_bits_7_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_7_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_7_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_7_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_7_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_7_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_8_din = io_is_current_tier ? io_out_din[287:256] : io_in_bits_8_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_8_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_8_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_8_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_8_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_8_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_9_din = io_is_current_tier ? io_out_din[319:288] : io_in_bits_9_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_9_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_9_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_9_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_9_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_9_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_10_din = io_is_current_tier ? io_out_din[351:320] : io_in_bits_10_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_10_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_10_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_10_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_10_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_10_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_11_din = io_is_current_tier ? io_out_din[383:352] : io_in_bits_11_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_11_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_11_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_11_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_11_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_11_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_12_din = io_is_current_tier ? io_out_din[415:384] : io_in_bits_12_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_12_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_12_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_12_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_12_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_12_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_13_din = io_is_current_tier ? io_out_din[447:416] : io_in_bits_13_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_13_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_13_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_13_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_13_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_13_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_14_din = io_is_current_tier ? io_out_din[479:448] : io_in_bits_14_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_14_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_14_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_14_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_14_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_14_srst = reset; // @[BFS.scala 1144:32]
  assign collector_fifos_15_din = io_is_current_tier ? io_out_din[511:480] : io_in_bits_15_tdata; // @[BFS.scala 1140:22]
  assign collector_fifos_15_wr_en = io_is_current_tier ? io_out_wr_en : io_in_valid & io_in_bits_15_tkeep; // @[BFS.scala 1141:24]
  assign collector_fifos_15_rd_en = io_out_rd_en; // @[BFS.scala 1145:18]
  assign collector_fifos_15_clk = clock; // @[BFS.scala 1143:31]
  assign collector_fifos_15_srst = reset; // @[BFS.scala 1144:32]
endmodule
module multi_port_mc(
  input          clock,
  input          reset,
  input          io_cacheable_out_ready,
  output         io_cacheable_out_valid,
  output [511:0] io_cacheable_out_bits_tdata,
  output [15:0]  io_cacheable_out_bits_tkeep,
  output         io_cacheable_in_0_ready,
  input          io_cacheable_in_0_valid,
  input  [31:0]  io_cacheable_in_0_bits_tdata,
  output         io_cacheable_in_1_ready,
  input          io_cacheable_in_1_valid,
  input  [31:0]  io_cacheable_in_1_bits_tdata,
  output         io_cacheable_in_2_ready,
  input          io_cacheable_in_2_valid,
  input  [31:0]  io_cacheable_in_2_bits_tdata,
  output         io_cacheable_in_3_ready,
  input          io_cacheable_in_3_valid,
  input  [31:0]  io_cacheable_in_3_bits_tdata,
  output         io_cacheable_in_4_ready,
  input          io_cacheable_in_4_valid,
  input  [31:0]  io_cacheable_in_4_bits_tdata,
  output         io_cacheable_in_5_ready,
  input          io_cacheable_in_5_valid,
  input  [31:0]  io_cacheable_in_5_bits_tdata,
  output         io_cacheable_in_6_ready,
  input          io_cacheable_in_6_valid,
  input  [31:0]  io_cacheable_in_6_bits_tdata,
  output         io_cacheable_in_7_ready,
  input          io_cacheable_in_7_valid,
  input  [31:0]  io_cacheable_in_7_bits_tdata,
  output         io_cacheable_in_8_ready,
  input          io_cacheable_in_8_valid,
  input  [31:0]  io_cacheable_in_8_bits_tdata,
  output         io_cacheable_in_9_ready,
  input          io_cacheable_in_9_valid,
  input  [31:0]  io_cacheable_in_9_bits_tdata,
  output         io_cacheable_in_10_ready,
  input          io_cacheable_in_10_valid,
  input  [31:0]  io_cacheable_in_10_bits_tdata,
  output         io_cacheable_in_11_ready,
  input          io_cacheable_in_11_valid,
  input  [31:0]  io_cacheable_in_11_bits_tdata,
  output         io_cacheable_in_12_ready,
  input          io_cacheable_in_12_valid,
  input  [31:0]  io_cacheable_in_12_bits_tdata,
  output         io_cacheable_in_13_ready,
  input          io_cacheable_in_13_valid,
  input  [31:0]  io_cacheable_in_13_bits_tdata,
  output         io_cacheable_in_14_ready,
  input          io_cacheable_in_14_valid,
  input  [31:0]  io_cacheable_in_14_bits_tdata,
  output         io_cacheable_in_15_ready,
  input          io_cacheable_in_15_valid,
  input  [31:0]  io_cacheable_in_15_bits_tdata,
  input          io_ddr_out_0_aw_ready,
  output         io_ddr_out_0_aw_valid,
  output [63:0]  io_ddr_out_0_aw_bits_awaddr,
  input          io_ddr_out_0_ar_ready,
  output         io_ddr_out_0_ar_valid,
  output [63:0]  io_ddr_out_0_ar_bits_araddr,
  input          io_ddr_out_0_w_ready,
  output         io_ddr_out_0_w_valid,
  output [511:0] io_ddr_out_0_w_bits_wdata,
  output         io_ddr_out_0_w_bits_wlast,
  input          io_ddr_out_0_r_valid,
  input  [511:0] io_ddr_out_0_r_bits_rdata,
  input          io_ddr_out_0_r_bits_rlast,
  input  [63:0]  io_tiers_base_addr_0,
  input  [63:0]  io_tiers_base_addr_1,
  output [31:0]  io_unvisited_size,
  input          io_start,
  input          io_signal,
  input          io_end,
  output         io_signal_ack
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  tier_fifo_0_clock; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_reset; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_ready; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_valid; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_0_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_0_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_1_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_1_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_2_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_2_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_3_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_3_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_4_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_4_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_5_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_5_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_6_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_6_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_7_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_7_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_8_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_8_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_9_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_9_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_10_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_10_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_11_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_11_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_12_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_12_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_13_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_13_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_14_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_14_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_0_io_in_bits_15_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_in_bits_15_tkeep; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_out_almost_full; // @[BFS.scala 1187:46]
  wire [511:0] tier_fifo_0_io_out_din; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_out_wr_en; // @[BFS.scala 1187:46]
  wire [511:0] tier_fifo_0_io_out_dout; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_out_rd_en; // @[BFS.scala 1187:46]
  wire [13:0] tier_fifo_0_io_out_data_count; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_out_valid; // @[BFS.scala 1187:46]
  wire  tier_fifo_0_io_is_current_tier; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_clock; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_reset; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_ready; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_valid; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_0_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_0_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_1_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_1_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_2_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_2_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_3_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_3_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_4_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_4_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_5_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_5_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_6_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_6_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_7_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_7_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_8_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_8_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_9_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_9_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_10_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_10_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_11_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_11_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_12_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_12_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_13_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_13_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_14_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_14_tkeep; // @[BFS.scala 1187:46]
  wire [31:0] tier_fifo_1_io_in_bits_15_tdata; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_in_bits_15_tkeep; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_out_almost_full; // @[BFS.scala 1187:46]
  wire [511:0] tier_fifo_1_io_out_din; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_out_wr_en; // @[BFS.scala 1187:46]
  wire [511:0] tier_fifo_1_io_out_dout; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_out_rd_en; // @[BFS.scala 1187:46]
  wire [13:0] tier_fifo_1_io_out_data_count; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_out_valid; // @[BFS.scala 1187:46]
  wire  tier_fifo_1_io_is_current_tier; // @[BFS.scala 1187:46]
  wire  in_pipeline_0_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_0_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_0_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_0_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_0_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_0_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_0_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_0_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_0_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_0_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_0_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_0_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_1_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_1_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_1_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_1_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_1_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_1_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_1_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_1_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_1_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_1_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_1_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_1_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_2_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_2_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_2_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_2_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_2_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_2_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_2_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_2_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_2_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_2_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_2_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_2_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_3_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_3_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_3_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_3_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_3_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_3_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_3_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_3_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_3_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_3_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_3_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_3_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_4_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_4_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_4_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_4_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_4_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_4_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_4_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_4_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_4_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_4_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_4_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_4_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_5_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_5_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_5_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_5_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_5_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_5_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_5_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_5_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_5_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_5_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_5_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_5_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_6_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_6_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_6_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_6_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_6_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_6_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_6_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_6_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_6_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_6_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_6_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_6_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_7_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_7_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_7_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_7_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_7_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_7_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_7_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_7_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_7_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_7_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_7_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_7_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_8_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_8_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_8_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_8_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_8_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_8_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_8_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_8_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_8_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_8_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_8_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_8_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_9_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_9_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_9_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_9_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_9_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_9_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_9_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_9_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_9_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_9_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_9_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_9_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_10_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_10_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_10_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_10_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_10_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_10_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_10_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_10_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_10_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_10_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_10_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_10_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_11_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_11_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_11_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_11_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_11_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_11_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_11_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_11_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_11_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_11_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_11_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_11_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_12_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_12_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_12_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_12_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_12_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_12_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_12_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_12_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_12_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_12_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_12_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_12_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_13_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_13_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_13_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_13_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_13_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_13_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_13_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_13_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_13_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_13_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_13_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_13_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_14_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_14_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_14_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_14_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_14_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_14_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_14_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_14_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_14_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_14_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_14_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_14_m_axis_tlast; // @[BFS.scala 1267:11]
  wire  in_pipeline_15_aclk; // @[BFS.scala 1267:11]
  wire  in_pipeline_15_aresetn; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_15_s_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_15_s_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_15_s_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_15_s_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_15_s_axis_tlast; // @[BFS.scala 1267:11]
  wire [31:0] in_pipeline_15_m_axis_tdata; // @[BFS.scala 1267:11]
  wire [3:0] in_pipeline_15_m_axis_tkeep; // @[BFS.scala 1267:11]
  wire  in_pipeline_15_m_axis_tvalid; // @[BFS.scala 1267:11]
  wire  in_pipeline_15_m_axis_tready; // @[BFS.scala 1267:11]
  wire  in_pipeline_15_m_axis_tlast; // @[BFS.scala 1267:11]
  reg [31:0] tier_counter_0; // @[BFS.scala 1188:29]
  reg [31:0] tier_counter_1; // @[BFS.scala 1188:29]
  reg [4:0] status; // @[BFS.scala 1206:23]
  reg [4:0] tier_status_0; // @[BFS.scala 1207:28]
  reg [4:0] tier_status_1; // @[BFS.scala 1207:28]
  wire  _T_1 = io_start & status == 5'h0; // @[BFS.scala 1209:17]
  wire  _T_2 = status == 5'h2; // @[BFS.scala 1211:21]
  wire  _T_5 = status == 5'h5; // @[BFS.scala 1213:21]
  wire  _T_8 = status == 5'h7; // @[BFS.scala 1215:34]
  wire [4:0] _GEN_0 = tier_status_1 != 5'h0 ? 5'h12 : 5'h1; // @[BFS.scala 1216:39 BFS.scala 1217:14 BFS.scala 1219:14]
  wire  _T_11 = status == 5'h1; // @[BFS.scala 1221:21]
  wire  _T_14 = status == 5'h6; // @[BFS.scala 1223:21]
  wire  _T_17 = status == 5'h8; // @[BFS.scala 1225:34]
  wire [4:0] _GEN_1 = tier_status_0 != 5'h0 ? 5'h11 : 5'h2; // @[BFS.scala 1226:38 BFS.scala 1227:14 BFS.scala 1229:14]
  wire  _T_20 = status == 5'h11; // @[BFS.scala 1231:21]
  wire  _T_21 = tier_status_0 == 5'h0; // @[BFS.scala 1231:60]
  wire  _T_23 = status == 5'h12; // @[BFS.scala 1233:21]
  wire  _T_24 = tier_status_1 == 5'h0; // @[BFS.scala 1233:60]
  wire [4:0] _GEN_2 = io_end ? 5'h0 : status; // @[BFS.scala 1235:21 BFS.scala 1236:12 BFS.scala 1206:23]
  wire [4:0] _GEN_3 = status == 5'h12 & tier_status_1 == 5'h0 ? 5'h1 : _GEN_2; // @[BFS.scala 1233:73 BFS.scala 1234:12]
  wire [4:0] _GEN_4 = status == 5'h11 & tier_status_0 == 5'h0 ? 5'h2 : _GEN_3; // @[BFS.scala 1231:73 BFS.scala 1232:12]
  wire [4:0] _GEN_5 = io_signal & status == 5'h8 ? _GEN_1 : _GEN_4; // @[BFS.scala 1225:55]
  wire [4:0] _GEN_6 = status == 5'h6 & io_cacheable_out_valid & io_cacheable_out_ready ? 5'h8 : _GEN_5; // @[BFS.scala 1223:92 BFS.scala 1224:12]
  wire [4:0] _GEN_7 = status == 5'h1 & tier_counter_1 == 32'h0 ? 5'h6 : _GEN_6; // @[BFS.scala 1221:70 BFS.scala 1222:12]
  wire [4:0] _GEN_8 = io_signal & status == 5'h7 ? _GEN_0 : _GEN_7; // @[BFS.scala 1215:55]
  wire  next_tier_mask_hi = _T_2 | _T_5 | _T_8 | _T_23; // @[BFS.scala 1239:115]
  wire  next_tier_mask_lo = _T_11 | _T_14 | _T_17 | _T_20; // @[BFS.scala 1240:94]
  wire [1:0] next_tier_mask = {next_tier_mask_hi,next_tier_mask_lo}; // @[Cat.scala 30:58]
  reg [63:0] tier_base_addr_0; // @[BFS.scala 1242:31]
  reg [63:0] tier_base_addr_1; // @[BFS.scala 1242:31]
  wire  step_fin = io_signal & (_T_8 | _T_17); // @[BFS.scala 1243:28]
  wire  _axi_aw_valid_T_1 = tier_status_0 == 5'h3; // @[BFS.scala 1370:57]
  wire  _axi_aw_valid_T_2 = tier_status_1 == 5'h3; // @[BFS.scala 1370:90]
  wire  axi_aw_valid = next_tier_mask[0] ? tier_status_0 == 5'h3 : tier_status_1 == 5'h3; // @[BFS.scala 1370:22]
  wire [63:0] _tier_base_addr_0_T_1 = tier_base_addr_0 + 64'h400; // @[BFS.scala 1249:16]
  wire  _T_35 = ~next_tier_mask[0]; // @[BFS.scala 1250:18]
  wire  _axi_ar_valid_T_1 = tier_status_1 == 5'h4; // @[BFS.scala 1377:57]
  wire  _axi_ar_valid_T_2 = tier_status_0 == 5'h4; // @[BFS.scala 1377:89]
  wire  axi_ar_valid = next_tier_mask[0] ? tier_status_1 == 5'h4 : tier_status_0 == 5'h4; // @[BFS.scala 1377:22]
  wire [63:0] _tier_base_addr_1_T_1 = tier_base_addr_1 + 64'h400; // @[BFS.scala 1249:16]
  wire  _T_49 = ~next_tier_mask[1]; // @[BFS.scala 1250:18]
  wire  _T_55 = io_cacheable_in_0_ready & io_cacheable_in_0_valid; // @[BFS.scala 1257:72]
  wire  _T_56 = io_cacheable_in_1_ready & io_cacheable_in_1_valid; // @[BFS.scala 1257:72]
  wire  _T_57 = io_cacheable_in_2_ready & io_cacheable_in_2_valid; // @[BFS.scala 1257:72]
  wire  _T_58 = io_cacheable_in_3_ready & io_cacheable_in_3_valid; // @[BFS.scala 1257:72]
  wire  _T_59 = io_cacheable_in_4_ready & io_cacheable_in_4_valid; // @[BFS.scala 1257:72]
  wire  _T_60 = io_cacheable_in_5_ready & io_cacheable_in_5_valid; // @[BFS.scala 1257:72]
  wire  _T_61 = io_cacheable_in_6_ready & io_cacheable_in_6_valid; // @[BFS.scala 1257:72]
  wire  _T_62 = io_cacheable_in_7_ready & io_cacheable_in_7_valid; // @[BFS.scala 1257:72]
  wire  _T_63 = io_cacheable_in_8_ready & io_cacheable_in_8_valid; // @[BFS.scala 1257:72]
  wire  _T_64 = io_cacheable_in_9_ready & io_cacheable_in_9_valid; // @[BFS.scala 1257:72]
  wire  _T_65 = io_cacheable_in_10_ready & io_cacheable_in_10_valid; // @[BFS.scala 1257:72]
  wire  _T_66 = io_cacheable_in_11_ready & io_cacheable_in_11_valid; // @[BFS.scala 1257:72]
  wire  _T_67 = io_cacheable_in_12_ready & io_cacheable_in_12_valid; // @[BFS.scala 1257:72]
  wire  _T_68 = io_cacheable_in_13_ready & io_cacheable_in_13_valid; // @[BFS.scala 1257:72]
  wire  _T_69 = io_cacheable_in_14_ready & io_cacheable_in_14_valid; // @[BFS.scala 1257:72]
  wire  _T_70 = io_cacheable_in_15_ready & io_cacheable_in_15_valid; // @[BFS.scala 1257:72]
  wire  _T_85 = io_cacheable_in_0_ready & io_cacheable_in_0_valid | io_cacheable_in_1_ready & io_cacheable_in_1_valid |
    io_cacheable_in_2_ready & io_cacheable_in_2_valid | io_cacheable_in_3_ready & io_cacheable_in_3_valid |
    io_cacheable_in_4_ready & io_cacheable_in_4_valid | io_cacheable_in_5_ready & io_cacheable_in_5_valid |
    io_cacheable_in_6_ready & io_cacheable_in_6_valid | io_cacheable_in_7_ready & io_cacheable_in_7_valid |
    io_cacheable_in_8_ready & io_cacheable_in_8_valid | io_cacheable_in_9_ready & io_cacheable_in_9_valid |
    io_cacheable_in_10_ready & io_cacheable_in_10_valid | io_cacheable_in_11_ready & io_cacheable_in_11_valid |
    io_cacheable_in_12_ready & io_cacheable_in_12_valid | io_cacheable_in_13_ready & io_cacheable_in_13_valid |
    io_cacheable_in_14_ready & io_cacheable_in_14_valid | _T_70; // @[BFS.scala 1257:93]
  wire [5:0] _tier_counter_0_WIRE = {{5'd0}, _T_55}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_WIRE_1 = {{5'd0}, _T_56}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_17 = _tier_counter_0_WIRE + _tier_counter_0_WIRE_1; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_2 = {{5'd0}, _T_57}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_19 = _tier_counter_0_T_17 + _tier_counter_0_WIRE_2; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_3 = {{5'd0}, _T_58}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_21 = _tier_counter_0_T_19 + _tier_counter_0_WIRE_3; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_4 = {{5'd0}, _T_59}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_23 = _tier_counter_0_T_21 + _tier_counter_0_WIRE_4; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_5 = {{5'd0}, _T_60}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_25 = _tier_counter_0_T_23 + _tier_counter_0_WIRE_5; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_6 = {{5'd0}, _T_61}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_27 = _tier_counter_0_T_25 + _tier_counter_0_WIRE_6; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_7 = {{5'd0}, _T_62}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_29 = _tier_counter_0_T_27 + _tier_counter_0_WIRE_7; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_8 = {{5'd0}, _T_63}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_31 = _tier_counter_0_T_29 + _tier_counter_0_WIRE_8; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_9 = {{5'd0}, _T_64}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_33 = _tier_counter_0_T_31 + _tier_counter_0_WIRE_9; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_10 = {{5'd0}, _T_65}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_35 = _tier_counter_0_T_33 + _tier_counter_0_WIRE_10; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_11 = {{5'd0}, _T_66}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_37 = _tier_counter_0_T_35 + _tier_counter_0_WIRE_11; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_12 = {{5'd0}, _T_67}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_39 = _tier_counter_0_T_37 + _tier_counter_0_WIRE_12; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_13 = {{5'd0}, _T_68}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_41 = _tier_counter_0_T_39 + _tier_counter_0_WIRE_13; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_14 = {{5'd0}, _T_69}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_43 = _tier_counter_0_T_41 + _tier_counter_0_WIRE_14; // @[BFS.scala 1258:100]
  wire [5:0] _tier_counter_0_WIRE_15 = {{5'd0}, _T_70}; // @[BFS.scala 1258:78 BFS.scala 1258:78]
  wire [5:0] _tier_counter_0_T_45 = _tier_counter_0_T_43 + _tier_counter_0_WIRE_15; // @[BFS.scala 1258:100]
  wire [31:0] _GEN_39 = {{26'd0}, _tier_counter_0_T_45}; // @[BFS.scala 1258:16]
  wire [31:0] _tier_counter_0_T_47 = tier_counter_0 + _GEN_39; // @[BFS.scala 1258:16]
  wire [31:0] _tier_counter_0_T_50 = tier_counter_0 - 32'h10; // @[BFS.scala 1260:59]
  wire [31:0] _GEN_40 = {{18'd0}, tier_fifo_0_io_out_data_count}; // @[BFS.scala 1260:69]
  wire [31:0] _tier_counter_0_T_52 = tier_counter_0 - _GEN_40; // @[BFS.scala 1260:69]
  wire [31:0] _tier_counter_1_T_47 = tier_counter_1 + _GEN_39; // @[BFS.scala 1258:16]
  wire [31:0] _tier_counter_1_T_50 = tier_counter_1 - 32'h10; // @[BFS.scala 1260:59]
  wire [31:0] _GEN_42 = {{18'd0}, tier_fifo_1_io_out_data_count}; // @[BFS.scala 1260:69]
  wire [31:0] _tier_counter_1_T_52 = tier_counter_1 - _GEN_42; // @[BFS.scala 1260:69]
  wire  fifos_ready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  wire  _steps_T = in_pipeline_0_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_1 = in_pipeline_0_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire  _steps_T_4 = in_pipeline_1_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_5 = in_pipeline_1_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE = {{4'd0}, _steps_T_1}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] _steps_WIRE_1 = {{4'd0}, _steps_T_5}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_1 = _steps_WIRE + _steps_WIRE_1; // @[BFS.scala 1283:119]
  wire  _steps_T_11 = in_pipeline_2_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_12 = in_pipeline_2_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_4 = {{4'd0}, _steps_T_12}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_2 = steps_1 + _steps_WIRE_4; // @[BFS.scala 1283:119]
  wire  _steps_T_22 = in_pipeline_3_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_23 = in_pipeline_3_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_8 = {{4'd0}, _steps_T_23}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_3 = steps_2 + _steps_WIRE_8; // @[BFS.scala 1283:119]
  wire  _steps_T_37 = in_pipeline_4_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_38 = in_pipeline_4_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_13 = {{4'd0}, _steps_T_38}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_4 = steps_3 + _steps_WIRE_13; // @[BFS.scala 1283:119]
  wire  _steps_T_56 = in_pipeline_5_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_57 = in_pipeline_5_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_19 = {{4'd0}, _steps_T_57}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_5 = steps_4 + _steps_WIRE_19; // @[BFS.scala 1283:119]
  wire  _steps_T_79 = in_pipeline_6_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_80 = in_pipeline_6_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_26 = {{4'd0}, _steps_T_80}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_6 = steps_5 + _steps_WIRE_26; // @[BFS.scala 1283:119]
  wire  _steps_T_106 = in_pipeline_7_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_107 = in_pipeline_7_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_34 = {{4'd0}, _steps_T_107}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_7 = steps_6 + _steps_WIRE_34; // @[BFS.scala 1283:119]
  wire  _steps_T_137 = in_pipeline_8_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_138 = in_pipeline_8_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_43 = {{4'd0}, _steps_T_138}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_8 = steps_7 + _steps_WIRE_43; // @[BFS.scala 1283:119]
  wire  _steps_T_172 = in_pipeline_9_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_173 = in_pipeline_9_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_53 = {{4'd0}, _steps_T_173}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_9 = steps_8 + _steps_WIRE_53; // @[BFS.scala 1283:119]
  wire  _steps_T_211 = in_pipeline_10_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_212 = in_pipeline_10_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_64 = {{4'd0}, _steps_T_212}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_10 = steps_9 + _steps_WIRE_64; // @[BFS.scala 1283:119]
  wire  _steps_T_254 = in_pipeline_11_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_255 = in_pipeline_11_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_76 = {{4'd0}, _steps_T_255}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_11 = steps_10 + _steps_WIRE_76; // @[BFS.scala 1283:119]
  wire  _steps_T_301 = in_pipeline_12_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_302 = in_pipeline_12_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_89 = {{4'd0}, _steps_T_302}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_12 = steps_11 + _steps_WIRE_89; // @[BFS.scala 1283:119]
  wire  _steps_T_352 = in_pipeline_13_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_353 = in_pipeline_13_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_103 = {{4'd0}, _steps_T_353}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_13 = steps_12 + _steps_WIRE_103; // @[BFS.scala 1283:119]
  wire  _steps_T_407 = in_pipeline_14_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_408 = in_pipeline_14_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_118 = {{4'd0}, _steps_T_408}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_14 = steps_13 + _steps_WIRE_118; // @[BFS.scala 1283:119]
  wire  _steps_T_466 = in_pipeline_15_m_axis_tvalid; // @[BFS.scala 1283:71]
  wire  _steps_T_467 = in_pipeline_15_m_axis_tvalid & fifos_ready; // @[BFS.scala 1283:74]
  wire [4:0] _steps_WIRE_134 = {{4'd0}, _steps_T_467}; // @[BFS.scala 1283:98 BFS.scala 1283:98]
  wire [4:0] steps_15 = steps_14 + _steps_WIRE_134; // @[BFS.scala 1283:119]
  reg [9:0] counter; // @[BFS.scala 1286:24]
  wire [9:0] _GEN_43 = {{5'd0}, steps_15}; // @[BFS.scala 1181:15]
  wire [9:0] _counter_T_1 = counter + _GEN_43; // @[BFS.scala 1181:15]
  wire [9:0] _counter_T_6 = _counter_T_1 - 10'h10; // @[BFS.scala 1181:44]
  wire [9:0] _fifo_in_data_T_2 = 10'h0 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_4 = 10'h10 - counter; // @[BFS.scala 1184:49]
  wire [10:0] _fifo_in_data_T_5 = {{1'd0}, _fifo_in_data_T_4}; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_7 = counter <= 10'h0 ? _fifo_in_data_T_2 : _fifo_in_data_T_5[9:0]; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_9 = _fifo_in_data_T_7 + 10'h1; // @[BFS.scala 1294:39]
  wire [9:0] _GEN_46 = {{5'd0}, _steps_WIRE}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_10 = _fifo_in_data_T_9 == _GEN_46; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_47 = {{5'd0}, steps_1}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_21 = _fifo_in_data_T_9 == _GEN_47; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_48 = {{5'd0}, steps_2}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_32 = _fifo_in_data_T_9 == _GEN_48; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_49 = {{5'd0}, steps_3}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_43 = _fifo_in_data_T_9 == _GEN_49; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_50 = {{5'd0}, steps_4}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_54 = _fifo_in_data_T_9 == _GEN_50; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_51 = {{5'd0}, steps_5}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_65 = _fifo_in_data_T_9 == _GEN_51; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_52 = {{5'd0}, steps_6}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_76 = _fifo_in_data_T_9 == _GEN_52; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_53 = {{5'd0}, steps_7}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_87 = _fifo_in_data_T_9 == _GEN_53; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_54 = {{5'd0}, steps_8}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_98 = _fifo_in_data_T_9 == _GEN_54; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_55 = {{5'd0}, steps_9}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_109 = _fifo_in_data_T_9 == _GEN_55; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_56 = {{5'd0}, steps_10}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_120 = _fifo_in_data_T_9 == _GEN_56; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_57 = {{5'd0}, steps_11}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_131 = _fifo_in_data_T_9 == _GEN_57; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_58 = {{5'd0}, steps_12}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_142 = _fifo_in_data_T_9 == _GEN_58; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_59 = {{5'd0}, steps_13}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_153 = _fifo_in_data_T_9 == _GEN_59; // @[BFS.scala 1294:46]
  wire [9:0] _GEN_60 = {{5'd0}, steps_14}; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_164 = _fifo_in_data_T_9 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_175 = _fifo_in_data_T_9 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_176 = _fifo_in_data_T_175 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_177 = _fifo_in_data_T_164 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_176; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_178 = _fifo_in_data_T_153 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_177; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_179 = _fifo_in_data_T_142 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_178; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_180 = _fifo_in_data_T_131 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_179; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_181 = _fifo_in_data_T_120 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_180; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_182 = _fifo_in_data_T_109 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_181; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_183 = _fifo_in_data_T_98 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_182; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_184 = _fifo_in_data_T_87 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_183; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_185 = _fifo_in_data_T_76 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_184; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_186 = _fifo_in_data_T_65 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_185; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_187 = _fifo_in_data_T_54 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_186; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_188 = _fifo_in_data_T_43 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_187; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_189 = _fifo_in_data_T_32 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_188; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_190 = _fifo_in_data_T_21 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_189; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_193 = 10'h1 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_197 = _fifo_in_data_T_4 + 10'h1; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_198 = counter <= 10'h1 ? _fifo_in_data_T_193 : _fifo_in_data_T_197; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_200 = _fifo_in_data_T_198 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_201 = _fifo_in_data_T_200 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_212 = _fifo_in_data_T_200 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_223 = _fifo_in_data_T_200 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_234 = _fifo_in_data_T_200 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_245 = _fifo_in_data_T_200 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_256 = _fifo_in_data_T_200 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_267 = _fifo_in_data_T_200 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_278 = _fifo_in_data_T_200 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_289 = _fifo_in_data_T_200 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_300 = _fifo_in_data_T_200 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_311 = _fifo_in_data_T_200 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_322 = _fifo_in_data_T_200 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_333 = _fifo_in_data_T_200 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_344 = _fifo_in_data_T_200 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_355 = _fifo_in_data_T_200 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_366 = _fifo_in_data_T_200 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_367 = _fifo_in_data_T_366 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_368 = _fifo_in_data_T_355 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_367; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_369 = _fifo_in_data_T_344 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_368; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_370 = _fifo_in_data_T_333 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_369; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_371 = _fifo_in_data_T_322 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_370; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_372 = _fifo_in_data_T_311 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_371; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_373 = _fifo_in_data_T_300 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_372; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_374 = _fifo_in_data_T_289 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_373; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_375 = _fifo_in_data_T_278 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_374; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_376 = _fifo_in_data_T_267 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_375; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_377 = _fifo_in_data_T_256 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_376; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_378 = _fifo_in_data_T_245 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_377; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_379 = _fifo_in_data_T_234 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_378; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_380 = _fifo_in_data_T_223 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_379; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_381 = _fifo_in_data_T_212 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_380; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_384 = 10'h2 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_388 = _fifo_in_data_T_4 + 10'h2; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_389 = counter <= 10'h2 ? _fifo_in_data_T_384 : _fifo_in_data_T_388; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_391 = _fifo_in_data_T_389 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_392 = _fifo_in_data_T_391 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_403 = _fifo_in_data_T_391 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_414 = _fifo_in_data_T_391 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_425 = _fifo_in_data_T_391 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_436 = _fifo_in_data_T_391 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_447 = _fifo_in_data_T_391 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_458 = _fifo_in_data_T_391 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_469 = _fifo_in_data_T_391 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_480 = _fifo_in_data_T_391 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_491 = _fifo_in_data_T_391 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_502 = _fifo_in_data_T_391 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_513 = _fifo_in_data_T_391 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_524 = _fifo_in_data_T_391 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_535 = _fifo_in_data_T_391 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_546 = _fifo_in_data_T_391 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_557 = _fifo_in_data_T_391 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_558 = _fifo_in_data_T_557 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_559 = _fifo_in_data_T_546 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_558; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_560 = _fifo_in_data_T_535 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_559; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_561 = _fifo_in_data_T_524 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_560; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_562 = _fifo_in_data_T_513 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_561; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_563 = _fifo_in_data_T_502 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_562; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_564 = _fifo_in_data_T_491 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_563; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_565 = _fifo_in_data_T_480 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_564; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_566 = _fifo_in_data_T_469 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_565; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_567 = _fifo_in_data_T_458 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_566; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_568 = _fifo_in_data_T_447 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_567; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_569 = _fifo_in_data_T_436 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_568; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_570 = _fifo_in_data_T_425 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_569; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_571 = _fifo_in_data_T_414 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_570; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_572 = _fifo_in_data_T_403 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_571; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_575 = 10'h3 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_579 = _fifo_in_data_T_4 + 10'h3; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_580 = counter <= 10'h3 ? _fifo_in_data_T_575 : _fifo_in_data_T_579; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_582 = _fifo_in_data_T_580 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_583 = _fifo_in_data_T_582 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_594 = _fifo_in_data_T_582 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_605 = _fifo_in_data_T_582 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_616 = _fifo_in_data_T_582 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_627 = _fifo_in_data_T_582 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_638 = _fifo_in_data_T_582 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_649 = _fifo_in_data_T_582 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_660 = _fifo_in_data_T_582 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_671 = _fifo_in_data_T_582 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_682 = _fifo_in_data_T_582 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_693 = _fifo_in_data_T_582 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_704 = _fifo_in_data_T_582 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_715 = _fifo_in_data_T_582 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_726 = _fifo_in_data_T_582 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_737 = _fifo_in_data_T_582 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_748 = _fifo_in_data_T_582 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_749 = _fifo_in_data_T_748 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_750 = _fifo_in_data_T_737 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_749; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_751 = _fifo_in_data_T_726 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_750; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_752 = _fifo_in_data_T_715 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_751; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_753 = _fifo_in_data_T_704 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_752; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_754 = _fifo_in_data_T_693 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_753; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_755 = _fifo_in_data_T_682 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_754; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_756 = _fifo_in_data_T_671 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_755; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_757 = _fifo_in_data_T_660 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_756; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_758 = _fifo_in_data_T_649 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_757; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_759 = _fifo_in_data_T_638 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_758; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_760 = _fifo_in_data_T_627 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_759; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_761 = _fifo_in_data_T_616 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_760; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_762 = _fifo_in_data_T_605 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_761; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_763 = _fifo_in_data_T_594 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_762; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_766 = 10'h4 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_770 = _fifo_in_data_T_4 + 10'h4; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_771 = counter <= 10'h4 ? _fifo_in_data_T_766 : _fifo_in_data_T_770; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_773 = _fifo_in_data_T_771 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_774 = _fifo_in_data_T_773 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_785 = _fifo_in_data_T_773 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_796 = _fifo_in_data_T_773 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_807 = _fifo_in_data_T_773 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_818 = _fifo_in_data_T_773 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_829 = _fifo_in_data_T_773 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_840 = _fifo_in_data_T_773 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_851 = _fifo_in_data_T_773 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_862 = _fifo_in_data_T_773 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_873 = _fifo_in_data_T_773 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_884 = _fifo_in_data_T_773 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_895 = _fifo_in_data_T_773 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_906 = _fifo_in_data_T_773 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_917 = _fifo_in_data_T_773 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_928 = _fifo_in_data_T_773 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_939 = _fifo_in_data_T_773 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_940 = _fifo_in_data_T_939 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_941 = _fifo_in_data_T_928 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_940; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_942 = _fifo_in_data_T_917 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_941; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_943 = _fifo_in_data_T_906 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_942; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_944 = _fifo_in_data_T_895 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_943; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_945 = _fifo_in_data_T_884 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_944; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_946 = _fifo_in_data_T_873 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_945; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_947 = _fifo_in_data_T_862 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_946; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_948 = _fifo_in_data_T_851 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_947; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_949 = _fifo_in_data_T_840 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_948; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_950 = _fifo_in_data_T_829 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_949; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_951 = _fifo_in_data_T_818 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_950; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_952 = _fifo_in_data_T_807 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_951; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_953 = _fifo_in_data_T_796 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_952; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_954 = _fifo_in_data_T_785 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_953; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_957 = 10'h5 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_961 = _fifo_in_data_T_4 + 10'h5; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_962 = counter <= 10'h5 ? _fifo_in_data_T_957 : _fifo_in_data_T_961; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_964 = _fifo_in_data_T_962 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_965 = _fifo_in_data_T_964 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_976 = _fifo_in_data_T_964 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_987 = _fifo_in_data_T_964 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_998 = _fifo_in_data_T_964 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1009 = _fifo_in_data_T_964 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1020 = _fifo_in_data_T_964 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1031 = _fifo_in_data_T_964 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1042 = _fifo_in_data_T_964 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1053 = _fifo_in_data_T_964 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1064 = _fifo_in_data_T_964 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1075 = _fifo_in_data_T_964 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1086 = _fifo_in_data_T_964 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1097 = _fifo_in_data_T_964 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1108 = _fifo_in_data_T_964 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1119 = _fifo_in_data_T_964 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1130 = _fifo_in_data_T_964 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_1131 = _fifo_in_data_T_1130 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1132 = _fifo_in_data_T_1119 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_1131; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1133 = _fifo_in_data_T_1108 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_1132; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1134 = _fifo_in_data_T_1097 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_1133; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1135 = _fifo_in_data_T_1086 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_1134; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1136 = _fifo_in_data_T_1075 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_1135; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1137 = _fifo_in_data_T_1064 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_1136; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1138 = _fifo_in_data_T_1053 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_1137; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1139 = _fifo_in_data_T_1042 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_1138; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1140 = _fifo_in_data_T_1031 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_1139; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1141 = _fifo_in_data_T_1020 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_1140; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1142 = _fifo_in_data_T_1009 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_1141; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1143 = _fifo_in_data_T_998 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_1142; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1144 = _fifo_in_data_T_987 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_1143; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1145 = _fifo_in_data_T_976 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_1144; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_1148 = 10'h6 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_1152 = _fifo_in_data_T_4 + 10'h6; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_1153 = counter <= 10'h6 ? _fifo_in_data_T_1148 : _fifo_in_data_T_1152; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_1155 = _fifo_in_data_T_1153 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_1156 = _fifo_in_data_T_1155 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1167 = _fifo_in_data_T_1155 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1178 = _fifo_in_data_T_1155 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1189 = _fifo_in_data_T_1155 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1200 = _fifo_in_data_T_1155 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1211 = _fifo_in_data_T_1155 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1222 = _fifo_in_data_T_1155 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1233 = _fifo_in_data_T_1155 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1244 = _fifo_in_data_T_1155 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1255 = _fifo_in_data_T_1155 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1266 = _fifo_in_data_T_1155 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1277 = _fifo_in_data_T_1155 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1288 = _fifo_in_data_T_1155 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1299 = _fifo_in_data_T_1155 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1310 = _fifo_in_data_T_1155 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1321 = _fifo_in_data_T_1155 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_1322 = _fifo_in_data_T_1321 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1323 = _fifo_in_data_T_1310 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_1322; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1324 = _fifo_in_data_T_1299 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_1323; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1325 = _fifo_in_data_T_1288 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_1324; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1326 = _fifo_in_data_T_1277 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_1325; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1327 = _fifo_in_data_T_1266 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_1326; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1328 = _fifo_in_data_T_1255 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_1327; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1329 = _fifo_in_data_T_1244 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_1328; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1330 = _fifo_in_data_T_1233 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_1329; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1331 = _fifo_in_data_T_1222 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_1330; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1332 = _fifo_in_data_T_1211 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_1331; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1333 = _fifo_in_data_T_1200 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_1332; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1334 = _fifo_in_data_T_1189 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_1333; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1335 = _fifo_in_data_T_1178 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_1334; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1336 = _fifo_in_data_T_1167 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_1335; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_1339 = 10'h7 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_1343 = _fifo_in_data_T_4 + 10'h7; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_1344 = counter <= 10'h7 ? _fifo_in_data_T_1339 : _fifo_in_data_T_1343; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_1346 = _fifo_in_data_T_1344 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_1347 = _fifo_in_data_T_1346 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1358 = _fifo_in_data_T_1346 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1369 = _fifo_in_data_T_1346 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1380 = _fifo_in_data_T_1346 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1391 = _fifo_in_data_T_1346 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1402 = _fifo_in_data_T_1346 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1413 = _fifo_in_data_T_1346 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1424 = _fifo_in_data_T_1346 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1435 = _fifo_in_data_T_1346 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1446 = _fifo_in_data_T_1346 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1457 = _fifo_in_data_T_1346 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1468 = _fifo_in_data_T_1346 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1479 = _fifo_in_data_T_1346 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1490 = _fifo_in_data_T_1346 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1501 = _fifo_in_data_T_1346 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1512 = _fifo_in_data_T_1346 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_1513 = _fifo_in_data_T_1512 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1514 = _fifo_in_data_T_1501 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_1513; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1515 = _fifo_in_data_T_1490 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_1514; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1516 = _fifo_in_data_T_1479 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_1515; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1517 = _fifo_in_data_T_1468 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_1516; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1518 = _fifo_in_data_T_1457 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_1517; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1519 = _fifo_in_data_T_1446 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_1518; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1520 = _fifo_in_data_T_1435 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_1519; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1521 = _fifo_in_data_T_1424 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_1520; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1522 = _fifo_in_data_T_1413 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_1521; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1523 = _fifo_in_data_T_1402 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_1522; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1524 = _fifo_in_data_T_1391 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_1523; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1525 = _fifo_in_data_T_1380 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_1524; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1526 = _fifo_in_data_T_1369 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_1525; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1527 = _fifo_in_data_T_1358 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_1526; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_1530 = 10'h8 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_1534 = _fifo_in_data_T_4 + 10'h8; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_1535 = counter <= 10'h8 ? _fifo_in_data_T_1530 : _fifo_in_data_T_1534; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_1537 = _fifo_in_data_T_1535 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_1538 = _fifo_in_data_T_1537 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1549 = _fifo_in_data_T_1537 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1560 = _fifo_in_data_T_1537 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1571 = _fifo_in_data_T_1537 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1582 = _fifo_in_data_T_1537 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1593 = _fifo_in_data_T_1537 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1604 = _fifo_in_data_T_1537 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1615 = _fifo_in_data_T_1537 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1626 = _fifo_in_data_T_1537 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1637 = _fifo_in_data_T_1537 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1648 = _fifo_in_data_T_1537 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1659 = _fifo_in_data_T_1537 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1670 = _fifo_in_data_T_1537 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1681 = _fifo_in_data_T_1537 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1692 = _fifo_in_data_T_1537 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1703 = _fifo_in_data_T_1537 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_1704 = _fifo_in_data_T_1703 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1705 = _fifo_in_data_T_1692 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_1704; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1706 = _fifo_in_data_T_1681 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_1705; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1707 = _fifo_in_data_T_1670 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_1706; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1708 = _fifo_in_data_T_1659 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_1707; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1709 = _fifo_in_data_T_1648 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_1708; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1710 = _fifo_in_data_T_1637 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_1709; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1711 = _fifo_in_data_T_1626 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_1710; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1712 = _fifo_in_data_T_1615 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_1711; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1713 = _fifo_in_data_T_1604 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_1712; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1714 = _fifo_in_data_T_1593 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_1713; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1715 = _fifo_in_data_T_1582 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_1714; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1716 = _fifo_in_data_T_1571 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_1715; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1717 = _fifo_in_data_T_1560 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_1716; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1718 = _fifo_in_data_T_1549 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_1717; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_1721 = 10'h9 - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_1725 = _fifo_in_data_T_4 + 10'h9; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_1726 = counter <= 10'h9 ? _fifo_in_data_T_1721 : _fifo_in_data_T_1725; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_1728 = _fifo_in_data_T_1726 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_1729 = _fifo_in_data_T_1728 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1740 = _fifo_in_data_T_1728 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1751 = _fifo_in_data_T_1728 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1762 = _fifo_in_data_T_1728 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1773 = _fifo_in_data_T_1728 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1784 = _fifo_in_data_T_1728 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1795 = _fifo_in_data_T_1728 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1806 = _fifo_in_data_T_1728 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1817 = _fifo_in_data_T_1728 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1828 = _fifo_in_data_T_1728 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1839 = _fifo_in_data_T_1728 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1850 = _fifo_in_data_T_1728 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1861 = _fifo_in_data_T_1728 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1872 = _fifo_in_data_T_1728 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1883 = _fifo_in_data_T_1728 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1894 = _fifo_in_data_T_1728 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_1895 = _fifo_in_data_T_1894 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1896 = _fifo_in_data_T_1883 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_1895; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1897 = _fifo_in_data_T_1872 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_1896; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1898 = _fifo_in_data_T_1861 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_1897; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1899 = _fifo_in_data_T_1850 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_1898; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1900 = _fifo_in_data_T_1839 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_1899; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1901 = _fifo_in_data_T_1828 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_1900; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1902 = _fifo_in_data_T_1817 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_1901; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1903 = _fifo_in_data_T_1806 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_1902; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1904 = _fifo_in_data_T_1795 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_1903; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1905 = _fifo_in_data_T_1784 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_1904; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1906 = _fifo_in_data_T_1773 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_1905; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1907 = _fifo_in_data_T_1762 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_1906; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1908 = _fifo_in_data_T_1751 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_1907; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1909 = _fifo_in_data_T_1740 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_1908; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_1912 = 10'ha - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_1916 = _fifo_in_data_T_4 + 10'ha; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_1917 = counter <= 10'ha ? _fifo_in_data_T_1912 : _fifo_in_data_T_1916; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_1919 = _fifo_in_data_T_1917 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_1920 = _fifo_in_data_T_1919 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1931 = _fifo_in_data_T_1919 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1942 = _fifo_in_data_T_1919 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1953 = _fifo_in_data_T_1919 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1964 = _fifo_in_data_T_1919 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1975 = _fifo_in_data_T_1919 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1986 = _fifo_in_data_T_1919 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_1997 = _fifo_in_data_T_1919 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2008 = _fifo_in_data_T_1919 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2019 = _fifo_in_data_T_1919 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2030 = _fifo_in_data_T_1919 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2041 = _fifo_in_data_T_1919 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2052 = _fifo_in_data_T_1919 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2063 = _fifo_in_data_T_1919 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2074 = _fifo_in_data_T_1919 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2085 = _fifo_in_data_T_1919 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_2086 = _fifo_in_data_T_2085 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2087 = _fifo_in_data_T_2074 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_2086; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2088 = _fifo_in_data_T_2063 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_2087; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2089 = _fifo_in_data_T_2052 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_2088; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2090 = _fifo_in_data_T_2041 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_2089; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2091 = _fifo_in_data_T_2030 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_2090; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2092 = _fifo_in_data_T_2019 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_2091; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2093 = _fifo_in_data_T_2008 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_2092; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2094 = _fifo_in_data_T_1997 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_2093; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2095 = _fifo_in_data_T_1986 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_2094; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2096 = _fifo_in_data_T_1975 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_2095; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2097 = _fifo_in_data_T_1964 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_2096; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2098 = _fifo_in_data_T_1953 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_2097; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2099 = _fifo_in_data_T_1942 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_2098; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2100 = _fifo_in_data_T_1931 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_2099; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_2103 = 10'hb - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_2107 = _fifo_in_data_T_4 + 10'hb; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_2108 = counter <= 10'hb ? _fifo_in_data_T_2103 : _fifo_in_data_T_2107; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_2110 = _fifo_in_data_T_2108 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_2111 = _fifo_in_data_T_2110 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2122 = _fifo_in_data_T_2110 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2133 = _fifo_in_data_T_2110 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2144 = _fifo_in_data_T_2110 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2155 = _fifo_in_data_T_2110 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2166 = _fifo_in_data_T_2110 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2177 = _fifo_in_data_T_2110 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2188 = _fifo_in_data_T_2110 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2199 = _fifo_in_data_T_2110 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2210 = _fifo_in_data_T_2110 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2221 = _fifo_in_data_T_2110 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2232 = _fifo_in_data_T_2110 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2243 = _fifo_in_data_T_2110 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2254 = _fifo_in_data_T_2110 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2265 = _fifo_in_data_T_2110 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2276 = _fifo_in_data_T_2110 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_2277 = _fifo_in_data_T_2276 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2278 = _fifo_in_data_T_2265 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_2277; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2279 = _fifo_in_data_T_2254 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_2278; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2280 = _fifo_in_data_T_2243 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_2279; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2281 = _fifo_in_data_T_2232 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_2280; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2282 = _fifo_in_data_T_2221 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_2281; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2283 = _fifo_in_data_T_2210 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_2282; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2284 = _fifo_in_data_T_2199 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_2283; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2285 = _fifo_in_data_T_2188 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_2284; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2286 = _fifo_in_data_T_2177 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_2285; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2287 = _fifo_in_data_T_2166 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_2286; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2288 = _fifo_in_data_T_2155 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_2287; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2289 = _fifo_in_data_T_2144 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_2288; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2290 = _fifo_in_data_T_2133 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_2289; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2291 = _fifo_in_data_T_2122 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_2290; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_2294 = 10'hc - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_2298 = _fifo_in_data_T_4 + 10'hc; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_2299 = counter <= 10'hc ? _fifo_in_data_T_2294 : _fifo_in_data_T_2298; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_2301 = _fifo_in_data_T_2299 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_2302 = _fifo_in_data_T_2301 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2313 = _fifo_in_data_T_2301 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2324 = _fifo_in_data_T_2301 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2335 = _fifo_in_data_T_2301 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2346 = _fifo_in_data_T_2301 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2357 = _fifo_in_data_T_2301 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2368 = _fifo_in_data_T_2301 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2379 = _fifo_in_data_T_2301 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2390 = _fifo_in_data_T_2301 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2401 = _fifo_in_data_T_2301 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2412 = _fifo_in_data_T_2301 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2423 = _fifo_in_data_T_2301 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2434 = _fifo_in_data_T_2301 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2445 = _fifo_in_data_T_2301 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2456 = _fifo_in_data_T_2301 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2467 = _fifo_in_data_T_2301 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_2468 = _fifo_in_data_T_2467 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2469 = _fifo_in_data_T_2456 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_2468; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2470 = _fifo_in_data_T_2445 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_2469; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2471 = _fifo_in_data_T_2434 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_2470; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2472 = _fifo_in_data_T_2423 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_2471; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2473 = _fifo_in_data_T_2412 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_2472; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2474 = _fifo_in_data_T_2401 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_2473; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2475 = _fifo_in_data_T_2390 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_2474; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2476 = _fifo_in_data_T_2379 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_2475; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2477 = _fifo_in_data_T_2368 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_2476; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2478 = _fifo_in_data_T_2357 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_2477; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2479 = _fifo_in_data_T_2346 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_2478; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2480 = _fifo_in_data_T_2335 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_2479; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2481 = _fifo_in_data_T_2324 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_2480; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2482 = _fifo_in_data_T_2313 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_2481; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_2485 = 10'hd - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_2489 = _fifo_in_data_T_4 + 10'hd; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_2490 = counter <= 10'hd ? _fifo_in_data_T_2485 : _fifo_in_data_T_2489; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_2492 = _fifo_in_data_T_2490 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_2493 = _fifo_in_data_T_2492 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2504 = _fifo_in_data_T_2492 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2515 = _fifo_in_data_T_2492 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2526 = _fifo_in_data_T_2492 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2537 = _fifo_in_data_T_2492 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2548 = _fifo_in_data_T_2492 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2559 = _fifo_in_data_T_2492 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2570 = _fifo_in_data_T_2492 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2581 = _fifo_in_data_T_2492 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2592 = _fifo_in_data_T_2492 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2603 = _fifo_in_data_T_2492 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2614 = _fifo_in_data_T_2492 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2625 = _fifo_in_data_T_2492 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2636 = _fifo_in_data_T_2492 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2647 = _fifo_in_data_T_2492 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2658 = _fifo_in_data_T_2492 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_2659 = _fifo_in_data_T_2658 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2660 = _fifo_in_data_T_2647 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_2659; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2661 = _fifo_in_data_T_2636 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_2660; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2662 = _fifo_in_data_T_2625 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_2661; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2663 = _fifo_in_data_T_2614 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_2662; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2664 = _fifo_in_data_T_2603 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_2663; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2665 = _fifo_in_data_T_2592 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_2664; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2666 = _fifo_in_data_T_2581 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_2665; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2667 = _fifo_in_data_T_2570 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_2666; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2668 = _fifo_in_data_T_2559 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_2667; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2669 = _fifo_in_data_T_2548 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_2668; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2670 = _fifo_in_data_T_2537 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_2669; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2671 = _fifo_in_data_T_2526 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_2670; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2672 = _fifo_in_data_T_2515 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_2671; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2673 = _fifo_in_data_T_2504 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_2672; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_2676 = 10'he - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_2680 = _fifo_in_data_T_4 + 10'he; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_2681 = counter <= 10'he ? _fifo_in_data_T_2676 : _fifo_in_data_T_2680; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_2683 = _fifo_in_data_T_2681 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_2684 = _fifo_in_data_T_2683 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2695 = _fifo_in_data_T_2683 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2706 = _fifo_in_data_T_2683 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2717 = _fifo_in_data_T_2683 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2728 = _fifo_in_data_T_2683 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2739 = _fifo_in_data_T_2683 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2750 = _fifo_in_data_T_2683 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2761 = _fifo_in_data_T_2683 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2772 = _fifo_in_data_T_2683 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2783 = _fifo_in_data_T_2683 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2794 = _fifo_in_data_T_2683 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2805 = _fifo_in_data_T_2683 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2816 = _fifo_in_data_T_2683 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2827 = _fifo_in_data_T_2683 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2838 = _fifo_in_data_T_2683 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2849 = _fifo_in_data_T_2683 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_2850 = _fifo_in_data_T_2849 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2851 = _fifo_in_data_T_2838 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_2850; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2852 = _fifo_in_data_T_2827 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_2851; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2853 = _fifo_in_data_T_2816 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_2852; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2854 = _fifo_in_data_T_2805 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_2853; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2855 = _fifo_in_data_T_2794 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_2854; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2856 = _fifo_in_data_T_2783 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_2855; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2857 = _fifo_in_data_T_2772 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_2856; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2858 = _fifo_in_data_T_2761 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_2857; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2859 = _fifo_in_data_T_2750 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_2858; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2860 = _fifo_in_data_T_2739 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_2859; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2861 = _fifo_in_data_T_2728 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_2860; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2862 = _fifo_in_data_T_2717 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_2861; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2863 = _fifo_in_data_T_2706 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_2862; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2864 = _fifo_in_data_T_2695 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_2863; // @[Mux.scala 98:16]
  wire [9:0] _fifo_in_data_T_2867 = 10'hf - counter; // @[BFS.scala 1184:34]
  wire [9:0] _fifo_in_data_T_2871 = _fifo_in_data_T_4 + 10'hf; // @[BFS.scala 1184:58]
  wire [9:0] _fifo_in_data_T_2872 = counter <= 10'hf ? _fifo_in_data_T_2867 : _fifo_in_data_T_2871; // @[BFS.scala 1184:8]
  wire [9:0] _fifo_in_data_T_2874 = _fifo_in_data_T_2872 + 10'h1; // @[BFS.scala 1294:39]
  wire  _fifo_in_data_T_2875 = _fifo_in_data_T_2874 == _GEN_46; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2886 = _fifo_in_data_T_2874 == _GEN_47; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2897 = _fifo_in_data_T_2874 == _GEN_48; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2908 = _fifo_in_data_T_2874 == _GEN_49; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2919 = _fifo_in_data_T_2874 == _GEN_50; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2930 = _fifo_in_data_T_2874 == _GEN_51; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2941 = _fifo_in_data_T_2874 == _GEN_52; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2952 = _fifo_in_data_T_2874 == _GEN_53; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2963 = _fifo_in_data_T_2874 == _GEN_54; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2974 = _fifo_in_data_T_2874 == _GEN_55; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2985 = _fifo_in_data_T_2874 == _GEN_56; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_2996 = _fifo_in_data_T_2874 == _GEN_57; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_3007 = _fifo_in_data_T_2874 == _GEN_58; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_3018 = _fifo_in_data_T_2874 == _GEN_59; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_3029 = _fifo_in_data_T_2874 == _GEN_60; // @[BFS.scala 1294:46]
  wire  _fifo_in_data_T_3040 = _fifo_in_data_T_2874 == _GEN_43; // @[BFS.scala 1294:46]
  wire [31:0] _fifo_in_data_T_3041 = _fifo_in_data_T_3040 ? in_pipeline_15_m_axis_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3042 = _fifo_in_data_T_3029 ? in_pipeline_14_m_axis_tdata : _fifo_in_data_T_3041; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3043 = _fifo_in_data_T_3018 ? in_pipeline_13_m_axis_tdata : _fifo_in_data_T_3042; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3044 = _fifo_in_data_T_3007 ? in_pipeline_12_m_axis_tdata : _fifo_in_data_T_3043; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3045 = _fifo_in_data_T_2996 ? in_pipeline_11_m_axis_tdata : _fifo_in_data_T_3044; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3046 = _fifo_in_data_T_2985 ? in_pipeline_10_m_axis_tdata : _fifo_in_data_T_3045; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3047 = _fifo_in_data_T_2974 ? in_pipeline_9_m_axis_tdata : _fifo_in_data_T_3046; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3048 = _fifo_in_data_T_2963 ? in_pipeline_8_m_axis_tdata : _fifo_in_data_T_3047; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3049 = _fifo_in_data_T_2952 ? in_pipeline_7_m_axis_tdata : _fifo_in_data_T_3048; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3050 = _fifo_in_data_T_2941 ? in_pipeline_6_m_axis_tdata : _fifo_in_data_T_3049; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3051 = _fifo_in_data_T_2930 ? in_pipeline_5_m_axis_tdata : _fifo_in_data_T_3050; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3052 = _fifo_in_data_T_2919 ? in_pipeline_4_m_axis_tdata : _fifo_in_data_T_3051; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3053 = _fifo_in_data_T_2908 ? in_pipeline_3_m_axis_tdata : _fifo_in_data_T_3052; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3054 = _fifo_in_data_T_2897 ? in_pipeline_2_m_axis_tdata : _fifo_in_data_T_3053; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3055 = _fifo_in_data_T_2886 ? in_pipeline_1_m_axis_tdata : _fifo_in_data_T_3054; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_193 = _fifo_in_data_T_164 ? _steps_T_407 : _fifo_in_data_T_175 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_194 = _fifo_in_data_T_153 ? _steps_T_352 : _fifo_in_valid_T_193; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_195 = _fifo_in_data_T_142 ? _steps_T_301 : _fifo_in_valid_T_194; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_196 = _fifo_in_data_T_131 ? _steps_T_254 : _fifo_in_valid_T_195; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_197 = _fifo_in_data_T_120 ? _steps_T_211 : _fifo_in_valid_T_196; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_198 = _fifo_in_data_T_109 ? _steps_T_172 : _fifo_in_valid_T_197; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_199 = _fifo_in_data_T_98 ? _steps_T_137 : _fifo_in_valid_T_198; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_200 = _fifo_in_data_T_87 ? _steps_T_106 : _fifo_in_valid_T_199; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_201 = _fifo_in_data_T_76 ? _steps_T_79 : _fifo_in_valid_T_200; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_202 = _fifo_in_data_T_65 ? _steps_T_56 : _fifo_in_valid_T_201; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_203 = _fifo_in_data_T_54 ? _steps_T_37 : _fifo_in_valid_T_202; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_204 = _fifo_in_data_T_43 ? _steps_T_22 : _fifo_in_valid_T_203; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_205 = _fifo_in_data_T_32 ? _steps_T_11 : _fifo_in_valid_T_204; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_206 = _fifo_in_data_T_21 ? _steps_T_4 : _fifo_in_valid_T_205; // @[Mux.scala 98:16]
  wire  fifo_in_valid_0 = _fifo_in_data_T_10 ? _steps_T : _fifo_in_valid_T_206; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_400 = _fifo_in_data_T_355 ? _steps_T_407 : _fifo_in_data_T_366 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_401 = _fifo_in_data_T_344 ? _steps_T_352 : _fifo_in_valid_T_400; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_402 = _fifo_in_data_T_333 ? _steps_T_301 : _fifo_in_valid_T_401; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_403 = _fifo_in_data_T_322 ? _steps_T_254 : _fifo_in_valid_T_402; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_404 = _fifo_in_data_T_311 ? _steps_T_211 : _fifo_in_valid_T_403; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_405 = _fifo_in_data_T_300 ? _steps_T_172 : _fifo_in_valid_T_404; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_406 = _fifo_in_data_T_289 ? _steps_T_137 : _fifo_in_valid_T_405; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_407 = _fifo_in_data_T_278 ? _steps_T_106 : _fifo_in_valid_T_406; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_408 = _fifo_in_data_T_267 ? _steps_T_79 : _fifo_in_valid_T_407; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_409 = _fifo_in_data_T_256 ? _steps_T_56 : _fifo_in_valid_T_408; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_410 = _fifo_in_data_T_245 ? _steps_T_37 : _fifo_in_valid_T_409; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_411 = _fifo_in_data_T_234 ? _steps_T_22 : _fifo_in_valid_T_410; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_412 = _fifo_in_data_T_223 ? _steps_T_11 : _fifo_in_valid_T_411; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_413 = _fifo_in_data_T_212 ? _steps_T_4 : _fifo_in_valid_T_412; // @[Mux.scala 98:16]
  wire  fifo_in_valid_1 = _fifo_in_data_T_201 ? _steps_T : _fifo_in_valid_T_413; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_607 = _fifo_in_data_T_546 ? _steps_T_407 : _fifo_in_data_T_557 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_608 = _fifo_in_data_T_535 ? _steps_T_352 : _fifo_in_valid_T_607; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_609 = _fifo_in_data_T_524 ? _steps_T_301 : _fifo_in_valid_T_608; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_610 = _fifo_in_data_T_513 ? _steps_T_254 : _fifo_in_valid_T_609; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_611 = _fifo_in_data_T_502 ? _steps_T_211 : _fifo_in_valid_T_610; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_612 = _fifo_in_data_T_491 ? _steps_T_172 : _fifo_in_valid_T_611; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_613 = _fifo_in_data_T_480 ? _steps_T_137 : _fifo_in_valid_T_612; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_614 = _fifo_in_data_T_469 ? _steps_T_106 : _fifo_in_valid_T_613; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_615 = _fifo_in_data_T_458 ? _steps_T_79 : _fifo_in_valid_T_614; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_616 = _fifo_in_data_T_447 ? _steps_T_56 : _fifo_in_valid_T_615; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_617 = _fifo_in_data_T_436 ? _steps_T_37 : _fifo_in_valid_T_616; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_618 = _fifo_in_data_T_425 ? _steps_T_22 : _fifo_in_valid_T_617; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_619 = _fifo_in_data_T_414 ? _steps_T_11 : _fifo_in_valid_T_618; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_620 = _fifo_in_data_T_403 ? _steps_T_4 : _fifo_in_valid_T_619; // @[Mux.scala 98:16]
  wire  fifo_in_valid_2 = _fifo_in_data_T_392 ? _steps_T : _fifo_in_valid_T_620; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_814 = _fifo_in_data_T_737 ? _steps_T_407 : _fifo_in_data_T_748 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_815 = _fifo_in_data_T_726 ? _steps_T_352 : _fifo_in_valid_T_814; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_816 = _fifo_in_data_T_715 ? _steps_T_301 : _fifo_in_valid_T_815; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_817 = _fifo_in_data_T_704 ? _steps_T_254 : _fifo_in_valid_T_816; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_818 = _fifo_in_data_T_693 ? _steps_T_211 : _fifo_in_valid_T_817; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_819 = _fifo_in_data_T_682 ? _steps_T_172 : _fifo_in_valid_T_818; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_820 = _fifo_in_data_T_671 ? _steps_T_137 : _fifo_in_valid_T_819; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_821 = _fifo_in_data_T_660 ? _steps_T_106 : _fifo_in_valid_T_820; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_822 = _fifo_in_data_T_649 ? _steps_T_79 : _fifo_in_valid_T_821; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_823 = _fifo_in_data_T_638 ? _steps_T_56 : _fifo_in_valid_T_822; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_824 = _fifo_in_data_T_627 ? _steps_T_37 : _fifo_in_valid_T_823; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_825 = _fifo_in_data_T_616 ? _steps_T_22 : _fifo_in_valid_T_824; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_826 = _fifo_in_data_T_605 ? _steps_T_11 : _fifo_in_valid_T_825; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_827 = _fifo_in_data_T_594 ? _steps_T_4 : _fifo_in_valid_T_826; // @[Mux.scala 98:16]
  wire  fifo_in_valid_3 = _fifo_in_data_T_583 ? _steps_T : _fifo_in_valid_T_827; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1021 = _fifo_in_data_T_928 ? _steps_T_407 : _fifo_in_data_T_939 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1022 = _fifo_in_data_T_917 ? _steps_T_352 : _fifo_in_valid_T_1021; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1023 = _fifo_in_data_T_906 ? _steps_T_301 : _fifo_in_valid_T_1022; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1024 = _fifo_in_data_T_895 ? _steps_T_254 : _fifo_in_valid_T_1023; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1025 = _fifo_in_data_T_884 ? _steps_T_211 : _fifo_in_valid_T_1024; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1026 = _fifo_in_data_T_873 ? _steps_T_172 : _fifo_in_valid_T_1025; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1027 = _fifo_in_data_T_862 ? _steps_T_137 : _fifo_in_valid_T_1026; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1028 = _fifo_in_data_T_851 ? _steps_T_106 : _fifo_in_valid_T_1027; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1029 = _fifo_in_data_T_840 ? _steps_T_79 : _fifo_in_valid_T_1028; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1030 = _fifo_in_data_T_829 ? _steps_T_56 : _fifo_in_valid_T_1029; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1031 = _fifo_in_data_T_818 ? _steps_T_37 : _fifo_in_valid_T_1030; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1032 = _fifo_in_data_T_807 ? _steps_T_22 : _fifo_in_valid_T_1031; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1033 = _fifo_in_data_T_796 ? _steps_T_11 : _fifo_in_valid_T_1032; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1034 = _fifo_in_data_T_785 ? _steps_T_4 : _fifo_in_valid_T_1033; // @[Mux.scala 98:16]
  wire  fifo_in_valid_4 = _fifo_in_data_T_774 ? _steps_T : _fifo_in_valid_T_1034; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1228 = _fifo_in_data_T_1119 ? _steps_T_407 : _fifo_in_data_T_1130 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1229 = _fifo_in_data_T_1108 ? _steps_T_352 : _fifo_in_valid_T_1228; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1230 = _fifo_in_data_T_1097 ? _steps_T_301 : _fifo_in_valid_T_1229; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1231 = _fifo_in_data_T_1086 ? _steps_T_254 : _fifo_in_valid_T_1230; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1232 = _fifo_in_data_T_1075 ? _steps_T_211 : _fifo_in_valid_T_1231; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1233 = _fifo_in_data_T_1064 ? _steps_T_172 : _fifo_in_valid_T_1232; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1234 = _fifo_in_data_T_1053 ? _steps_T_137 : _fifo_in_valid_T_1233; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1235 = _fifo_in_data_T_1042 ? _steps_T_106 : _fifo_in_valid_T_1234; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1236 = _fifo_in_data_T_1031 ? _steps_T_79 : _fifo_in_valid_T_1235; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1237 = _fifo_in_data_T_1020 ? _steps_T_56 : _fifo_in_valid_T_1236; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1238 = _fifo_in_data_T_1009 ? _steps_T_37 : _fifo_in_valid_T_1237; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1239 = _fifo_in_data_T_998 ? _steps_T_22 : _fifo_in_valid_T_1238; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1240 = _fifo_in_data_T_987 ? _steps_T_11 : _fifo_in_valid_T_1239; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1241 = _fifo_in_data_T_976 ? _steps_T_4 : _fifo_in_valid_T_1240; // @[Mux.scala 98:16]
  wire  fifo_in_valid_5 = _fifo_in_data_T_965 ? _steps_T : _fifo_in_valid_T_1241; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1435 = _fifo_in_data_T_1310 ? _steps_T_407 : _fifo_in_data_T_1321 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1436 = _fifo_in_data_T_1299 ? _steps_T_352 : _fifo_in_valid_T_1435; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1437 = _fifo_in_data_T_1288 ? _steps_T_301 : _fifo_in_valid_T_1436; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1438 = _fifo_in_data_T_1277 ? _steps_T_254 : _fifo_in_valid_T_1437; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1439 = _fifo_in_data_T_1266 ? _steps_T_211 : _fifo_in_valid_T_1438; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1440 = _fifo_in_data_T_1255 ? _steps_T_172 : _fifo_in_valid_T_1439; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1441 = _fifo_in_data_T_1244 ? _steps_T_137 : _fifo_in_valid_T_1440; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1442 = _fifo_in_data_T_1233 ? _steps_T_106 : _fifo_in_valid_T_1441; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1443 = _fifo_in_data_T_1222 ? _steps_T_79 : _fifo_in_valid_T_1442; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1444 = _fifo_in_data_T_1211 ? _steps_T_56 : _fifo_in_valid_T_1443; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1445 = _fifo_in_data_T_1200 ? _steps_T_37 : _fifo_in_valid_T_1444; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1446 = _fifo_in_data_T_1189 ? _steps_T_22 : _fifo_in_valid_T_1445; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1447 = _fifo_in_data_T_1178 ? _steps_T_11 : _fifo_in_valid_T_1446; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1448 = _fifo_in_data_T_1167 ? _steps_T_4 : _fifo_in_valid_T_1447; // @[Mux.scala 98:16]
  wire  fifo_in_valid_6 = _fifo_in_data_T_1156 ? _steps_T : _fifo_in_valid_T_1448; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1642 = _fifo_in_data_T_1501 ? _steps_T_407 : _fifo_in_data_T_1512 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1643 = _fifo_in_data_T_1490 ? _steps_T_352 : _fifo_in_valid_T_1642; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1644 = _fifo_in_data_T_1479 ? _steps_T_301 : _fifo_in_valid_T_1643; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1645 = _fifo_in_data_T_1468 ? _steps_T_254 : _fifo_in_valid_T_1644; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1646 = _fifo_in_data_T_1457 ? _steps_T_211 : _fifo_in_valid_T_1645; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1647 = _fifo_in_data_T_1446 ? _steps_T_172 : _fifo_in_valid_T_1646; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1648 = _fifo_in_data_T_1435 ? _steps_T_137 : _fifo_in_valid_T_1647; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1649 = _fifo_in_data_T_1424 ? _steps_T_106 : _fifo_in_valid_T_1648; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1650 = _fifo_in_data_T_1413 ? _steps_T_79 : _fifo_in_valid_T_1649; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1651 = _fifo_in_data_T_1402 ? _steps_T_56 : _fifo_in_valid_T_1650; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1652 = _fifo_in_data_T_1391 ? _steps_T_37 : _fifo_in_valid_T_1651; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1653 = _fifo_in_data_T_1380 ? _steps_T_22 : _fifo_in_valid_T_1652; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1654 = _fifo_in_data_T_1369 ? _steps_T_11 : _fifo_in_valid_T_1653; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1655 = _fifo_in_data_T_1358 ? _steps_T_4 : _fifo_in_valid_T_1654; // @[Mux.scala 98:16]
  wire  fifo_in_valid_7 = _fifo_in_data_T_1347 ? _steps_T : _fifo_in_valid_T_1655; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1849 = _fifo_in_data_T_1692 ? _steps_T_407 : _fifo_in_data_T_1703 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1850 = _fifo_in_data_T_1681 ? _steps_T_352 : _fifo_in_valid_T_1849; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1851 = _fifo_in_data_T_1670 ? _steps_T_301 : _fifo_in_valid_T_1850; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1852 = _fifo_in_data_T_1659 ? _steps_T_254 : _fifo_in_valid_T_1851; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1853 = _fifo_in_data_T_1648 ? _steps_T_211 : _fifo_in_valid_T_1852; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1854 = _fifo_in_data_T_1637 ? _steps_T_172 : _fifo_in_valid_T_1853; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1855 = _fifo_in_data_T_1626 ? _steps_T_137 : _fifo_in_valid_T_1854; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1856 = _fifo_in_data_T_1615 ? _steps_T_106 : _fifo_in_valid_T_1855; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1857 = _fifo_in_data_T_1604 ? _steps_T_79 : _fifo_in_valid_T_1856; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1858 = _fifo_in_data_T_1593 ? _steps_T_56 : _fifo_in_valid_T_1857; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1859 = _fifo_in_data_T_1582 ? _steps_T_37 : _fifo_in_valid_T_1858; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1860 = _fifo_in_data_T_1571 ? _steps_T_22 : _fifo_in_valid_T_1859; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1861 = _fifo_in_data_T_1560 ? _steps_T_11 : _fifo_in_valid_T_1860; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1862 = _fifo_in_data_T_1549 ? _steps_T_4 : _fifo_in_valid_T_1861; // @[Mux.scala 98:16]
  wire  fifo_in_valid_8 = _fifo_in_data_T_1538 ? _steps_T : _fifo_in_valid_T_1862; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2056 = _fifo_in_data_T_1883 ? _steps_T_407 : _fifo_in_data_T_1894 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2057 = _fifo_in_data_T_1872 ? _steps_T_352 : _fifo_in_valid_T_2056; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2058 = _fifo_in_data_T_1861 ? _steps_T_301 : _fifo_in_valid_T_2057; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2059 = _fifo_in_data_T_1850 ? _steps_T_254 : _fifo_in_valid_T_2058; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2060 = _fifo_in_data_T_1839 ? _steps_T_211 : _fifo_in_valid_T_2059; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2061 = _fifo_in_data_T_1828 ? _steps_T_172 : _fifo_in_valid_T_2060; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2062 = _fifo_in_data_T_1817 ? _steps_T_137 : _fifo_in_valid_T_2061; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2063 = _fifo_in_data_T_1806 ? _steps_T_106 : _fifo_in_valid_T_2062; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2064 = _fifo_in_data_T_1795 ? _steps_T_79 : _fifo_in_valid_T_2063; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2065 = _fifo_in_data_T_1784 ? _steps_T_56 : _fifo_in_valid_T_2064; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2066 = _fifo_in_data_T_1773 ? _steps_T_37 : _fifo_in_valid_T_2065; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2067 = _fifo_in_data_T_1762 ? _steps_T_22 : _fifo_in_valid_T_2066; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2068 = _fifo_in_data_T_1751 ? _steps_T_11 : _fifo_in_valid_T_2067; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2069 = _fifo_in_data_T_1740 ? _steps_T_4 : _fifo_in_valid_T_2068; // @[Mux.scala 98:16]
  wire  fifo_in_valid_9 = _fifo_in_data_T_1729 ? _steps_T : _fifo_in_valid_T_2069; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2263 = _fifo_in_data_T_2074 ? _steps_T_407 : _fifo_in_data_T_2085 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2264 = _fifo_in_data_T_2063 ? _steps_T_352 : _fifo_in_valid_T_2263; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2265 = _fifo_in_data_T_2052 ? _steps_T_301 : _fifo_in_valid_T_2264; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2266 = _fifo_in_data_T_2041 ? _steps_T_254 : _fifo_in_valid_T_2265; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2267 = _fifo_in_data_T_2030 ? _steps_T_211 : _fifo_in_valid_T_2266; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2268 = _fifo_in_data_T_2019 ? _steps_T_172 : _fifo_in_valid_T_2267; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2269 = _fifo_in_data_T_2008 ? _steps_T_137 : _fifo_in_valid_T_2268; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2270 = _fifo_in_data_T_1997 ? _steps_T_106 : _fifo_in_valid_T_2269; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2271 = _fifo_in_data_T_1986 ? _steps_T_79 : _fifo_in_valid_T_2270; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2272 = _fifo_in_data_T_1975 ? _steps_T_56 : _fifo_in_valid_T_2271; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2273 = _fifo_in_data_T_1964 ? _steps_T_37 : _fifo_in_valid_T_2272; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2274 = _fifo_in_data_T_1953 ? _steps_T_22 : _fifo_in_valid_T_2273; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2275 = _fifo_in_data_T_1942 ? _steps_T_11 : _fifo_in_valid_T_2274; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2276 = _fifo_in_data_T_1931 ? _steps_T_4 : _fifo_in_valid_T_2275; // @[Mux.scala 98:16]
  wire  fifo_in_valid_10 = _fifo_in_data_T_1920 ? _steps_T : _fifo_in_valid_T_2276; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2470 = _fifo_in_data_T_2265 ? _steps_T_407 : _fifo_in_data_T_2276 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2471 = _fifo_in_data_T_2254 ? _steps_T_352 : _fifo_in_valid_T_2470; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2472 = _fifo_in_data_T_2243 ? _steps_T_301 : _fifo_in_valid_T_2471; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2473 = _fifo_in_data_T_2232 ? _steps_T_254 : _fifo_in_valid_T_2472; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2474 = _fifo_in_data_T_2221 ? _steps_T_211 : _fifo_in_valid_T_2473; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2475 = _fifo_in_data_T_2210 ? _steps_T_172 : _fifo_in_valid_T_2474; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2476 = _fifo_in_data_T_2199 ? _steps_T_137 : _fifo_in_valid_T_2475; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2477 = _fifo_in_data_T_2188 ? _steps_T_106 : _fifo_in_valid_T_2476; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2478 = _fifo_in_data_T_2177 ? _steps_T_79 : _fifo_in_valid_T_2477; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2479 = _fifo_in_data_T_2166 ? _steps_T_56 : _fifo_in_valid_T_2478; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2480 = _fifo_in_data_T_2155 ? _steps_T_37 : _fifo_in_valid_T_2479; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2481 = _fifo_in_data_T_2144 ? _steps_T_22 : _fifo_in_valid_T_2480; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2482 = _fifo_in_data_T_2133 ? _steps_T_11 : _fifo_in_valid_T_2481; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2483 = _fifo_in_data_T_2122 ? _steps_T_4 : _fifo_in_valid_T_2482; // @[Mux.scala 98:16]
  wire  fifo_in_valid_11 = _fifo_in_data_T_2111 ? _steps_T : _fifo_in_valid_T_2483; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2677 = _fifo_in_data_T_2456 ? _steps_T_407 : _fifo_in_data_T_2467 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2678 = _fifo_in_data_T_2445 ? _steps_T_352 : _fifo_in_valid_T_2677; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2679 = _fifo_in_data_T_2434 ? _steps_T_301 : _fifo_in_valid_T_2678; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2680 = _fifo_in_data_T_2423 ? _steps_T_254 : _fifo_in_valid_T_2679; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2681 = _fifo_in_data_T_2412 ? _steps_T_211 : _fifo_in_valid_T_2680; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2682 = _fifo_in_data_T_2401 ? _steps_T_172 : _fifo_in_valid_T_2681; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2683 = _fifo_in_data_T_2390 ? _steps_T_137 : _fifo_in_valid_T_2682; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2684 = _fifo_in_data_T_2379 ? _steps_T_106 : _fifo_in_valid_T_2683; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2685 = _fifo_in_data_T_2368 ? _steps_T_79 : _fifo_in_valid_T_2684; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2686 = _fifo_in_data_T_2357 ? _steps_T_56 : _fifo_in_valid_T_2685; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2687 = _fifo_in_data_T_2346 ? _steps_T_37 : _fifo_in_valid_T_2686; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2688 = _fifo_in_data_T_2335 ? _steps_T_22 : _fifo_in_valid_T_2687; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2689 = _fifo_in_data_T_2324 ? _steps_T_11 : _fifo_in_valid_T_2688; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2690 = _fifo_in_data_T_2313 ? _steps_T_4 : _fifo_in_valid_T_2689; // @[Mux.scala 98:16]
  wire  fifo_in_valid_12 = _fifo_in_data_T_2302 ? _steps_T : _fifo_in_valid_T_2690; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2884 = _fifo_in_data_T_2647 ? _steps_T_407 : _fifo_in_data_T_2658 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2885 = _fifo_in_data_T_2636 ? _steps_T_352 : _fifo_in_valid_T_2884; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2886 = _fifo_in_data_T_2625 ? _steps_T_301 : _fifo_in_valid_T_2885; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2887 = _fifo_in_data_T_2614 ? _steps_T_254 : _fifo_in_valid_T_2886; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2888 = _fifo_in_data_T_2603 ? _steps_T_211 : _fifo_in_valid_T_2887; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2889 = _fifo_in_data_T_2592 ? _steps_T_172 : _fifo_in_valid_T_2888; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2890 = _fifo_in_data_T_2581 ? _steps_T_137 : _fifo_in_valid_T_2889; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2891 = _fifo_in_data_T_2570 ? _steps_T_106 : _fifo_in_valid_T_2890; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2892 = _fifo_in_data_T_2559 ? _steps_T_79 : _fifo_in_valid_T_2891; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2893 = _fifo_in_data_T_2548 ? _steps_T_56 : _fifo_in_valid_T_2892; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2894 = _fifo_in_data_T_2537 ? _steps_T_37 : _fifo_in_valid_T_2893; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2895 = _fifo_in_data_T_2526 ? _steps_T_22 : _fifo_in_valid_T_2894; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2896 = _fifo_in_data_T_2515 ? _steps_T_11 : _fifo_in_valid_T_2895; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2897 = _fifo_in_data_T_2504 ? _steps_T_4 : _fifo_in_valid_T_2896; // @[Mux.scala 98:16]
  wire  fifo_in_valid_13 = _fifo_in_data_T_2493 ? _steps_T : _fifo_in_valid_T_2897; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3091 = _fifo_in_data_T_2838 ? _steps_T_407 : _fifo_in_data_T_2849 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3092 = _fifo_in_data_T_2827 ? _steps_T_352 : _fifo_in_valid_T_3091; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3093 = _fifo_in_data_T_2816 ? _steps_T_301 : _fifo_in_valid_T_3092; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3094 = _fifo_in_data_T_2805 ? _steps_T_254 : _fifo_in_valid_T_3093; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3095 = _fifo_in_data_T_2794 ? _steps_T_211 : _fifo_in_valid_T_3094; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3096 = _fifo_in_data_T_2783 ? _steps_T_172 : _fifo_in_valid_T_3095; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3097 = _fifo_in_data_T_2772 ? _steps_T_137 : _fifo_in_valid_T_3096; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3098 = _fifo_in_data_T_2761 ? _steps_T_106 : _fifo_in_valid_T_3097; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3099 = _fifo_in_data_T_2750 ? _steps_T_79 : _fifo_in_valid_T_3098; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3100 = _fifo_in_data_T_2739 ? _steps_T_56 : _fifo_in_valid_T_3099; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3101 = _fifo_in_data_T_2728 ? _steps_T_37 : _fifo_in_valid_T_3100; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3102 = _fifo_in_data_T_2717 ? _steps_T_22 : _fifo_in_valid_T_3101; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3103 = _fifo_in_data_T_2706 ? _steps_T_11 : _fifo_in_valid_T_3102; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3104 = _fifo_in_data_T_2695 ? _steps_T_4 : _fifo_in_valid_T_3103; // @[Mux.scala 98:16]
  wire  fifo_in_valid_14 = _fifo_in_data_T_2684 ? _steps_T : _fifo_in_valid_T_3104; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3298 = _fifo_in_data_T_3029 ? _steps_T_407 : _fifo_in_data_T_3040 & _steps_T_466; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3299 = _fifo_in_data_T_3018 ? _steps_T_352 : _fifo_in_valid_T_3298; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3300 = _fifo_in_data_T_3007 ? _steps_T_301 : _fifo_in_valid_T_3299; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3301 = _fifo_in_data_T_2996 ? _steps_T_254 : _fifo_in_valid_T_3300; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3302 = _fifo_in_data_T_2985 ? _steps_T_211 : _fifo_in_valid_T_3301; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3303 = _fifo_in_data_T_2974 ? _steps_T_172 : _fifo_in_valid_T_3302; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3304 = _fifo_in_data_T_2963 ? _steps_T_137 : _fifo_in_valid_T_3303; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3305 = _fifo_in_data_T_2952 ? _steps_T_106 : _fifo_in_valid_T_3304; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3306 = _fifo_in_data_T_2941 ? _steps_T_79 : _fifo_in_valid_T_3305; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3307 = _fifo_in_data_T_2930 ? _steps_T_56 : _fifo_in_valid_T_3306; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3308 = _fifo_in_data_T_2919 ? _steps_T_37 : _fifo_in_valid_T_3307; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3309 = _fifo_in_data_T_2908 ? _steps_T_22 : _fifo_in_valid_T_3308; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3310 = _fifo_in_data_T_2897 ? _steps_T_11 : _fifo_in_valid_T_3309; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3311 = _fifo_in_data_T_2886 ? _steps_T_4 : _fifo_in_valid_T_3310; // @[Mux.scala 98:16]
  wire  fifo_in_valid_15 = _fifo_in_data_T_2875 ? _steps_T : _fifo_in_valid_T_3311; // @[Mux.scala 98:16]
    (*dont_touch = "true" *)reg [31:0] ready_counter; // @[BFS.scala 1302:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 1305:36]
  wire  _axi_w_valid_T_1 = tier_status_0 == 5'h9; // @[BFS.scala 1379:56]
  wire  _axi_w_valid_T_2 = tier_status_1 == 5'h9; // @[BFS.scala 1379:93]
  wire  axi_w_valid = next_tier_mask[0] ? tier_status_0 == 5'h9 : tier_status_1 == 5'h9; // @[BFS.scala 1379:21]
  wire  _tier_fifo_0_io_out_rd_en_T_3 = axi_w_valid & io_ddr_out_0_w_ready; // @[BFS.scala 1309:69]
  wire  _tier_fifo_0_io_out_rd_en_T_4 = io_cacheable_out_ready & io_cacheable_out_valid; // @[BFS.scala 1310:8]
  wire  _T_169 = next_tier_mask[0] & tier_fifo_0_io_out_almost_full & _T_21; // @[BFS.scala 1326:65]
  wire  _T_176 = tier_fifo_0_io_out_data_count == 14'h0; // @[BFS.scala 1126:23]
  reg [7:0] wcount; // @[BFS.scala 1358:23]
  wire  axi_w_bits_wlast = wcount == 8'h1; // @[BFS.scala 1380:30]
  wire [4:0] _GEN_25 = _axi_w_valid_T_1 & axi_w_bits_wlast & io_ddr_out_0_w_ready ? 5'h0 : tier_status_0; // @[BFS.scala 1337:94 BFS.scala 1338:11 BFS.scala 1207:28]
  wire [4:0] _GEN_26 = tier_status_0 == 5'h10 & io_ddr_out_0_r_bits_rlast & io_ddr_out_0_r_valid ? 5'h0 : _GEN_25; // @[BFS.scala 1335:99 BFS.scala 1336:11]
  wire [4:0] _GEN_27 = _axi_ar_valid_T_2 & io_ddr_out_0_ar_ready ? 5'h10 : _GEN_26; // @[BFS.scala 1333:52 BFS.scala 1334:11]
  wire  _T_199 = next_tier_mask[1] & tier_fifo_1_io_out_almost_full & _T_24; // @[BFS.scala 1326:65]
  wire  _T_206 = tier_fifo_1_io_out_data_count == 14'h0; // @[BFS.scala 1126:23]
  wire [4:0] _GEN_31 = _axi_w_valid_T_2 & axi_w_bits_wlast & io_ddr_out_0_w_ready ? 5'h0 : tier_status_1; // @[BFS.scala 1337:94 BFS.scala 1338:11 BFS.scala 1207:28]
  wire [4:0] _GEN_32 = tier_status_1 == 5'h10 & io_ddr_out_0_r_bits_rlast & io_ddr_out_0_r_valid ? 5'h0 : _GEN_31; // @[BFS.scala 1335:99 BFS.scala 1336:11]
  wire [4:0] _GEN_33 = _axi_ar_valid_T_1 & io_ddr_out_0_ar_ready ? 5'h10 : _GEN_32; // @[BFS.scala 1333:52 BFS.scala 1334:11]
  wire  _io_cacheable_out_valid_T_2 = tier_fifo_1_io_out_valid | _T_14; // @[BFS.scala 1345:57]
  wire  _io_cacheable_out_valid_T_5 = tier_fifo_0_io_out_valid | _T_5; // @[BFS.scala 1346:57]
  wire [511:0] _io_cacheable_out_bits_tdata_T_4 = next_tier_mask[1] ? tier_fifo_0_io_out_dout : 512'h0; // @[Mux.scala 98:16]
  wire [511:0] _io_cacheable_out_bits_tdata_T_5 = next_tier_mask[0] ? tier_fifo_1_io_out_dout :
    _io_cacheable_out_bits_tdata_T_4; // @[Mux.scala 98:16]
  wire [511:0] _io_cacheable_out_bits_tdata_T_6 = _T_14 ? 512'h80000000 : _io_cacheable_out_bits_tdata_T_5; // @[Mux.scala 98:16]
  wire  _io_cacheable_out_bits_tkeep_T_6 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h0 :
    tier_fifo_0_io_out_data_count > 14'h0; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_10 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h1 :
    tier_fifo_0_io_out_data_count > 14'h1; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_14 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h2 :
    tier_fifo_0_io_out_data_count > 14'h2; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_18 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h3 :
    tier_fifo_0_io_out_data_count > 14'h3; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_22 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h4 :
    tier_fifo_0_io_out_data_count > 14'h4; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_26 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h5 :
    tier_fifo_0_io_out_data_count > 14'h5; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_30 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h6 :
    tier_fifo_0_io_out_data_count > 14'h6; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_34 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h7 :
    tier_fifo_0_io_out_data_count > 14'h7; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_38 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h8 :
    tier_fifo_0_io_out_data_count > 14'h8; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_42 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'h9 :
    tier_fifo_0_io_out_data_count > 14'h9; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_46 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'ha :
    tier_fifo_0_io_out_data_count > 14'ha; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_50 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'hb :
    tier_fifo_0_io_out_data_count > 14'hb; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_54 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'hc :
    tier_fifo_0_io_out_data_count > 14'hc; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_58 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'hd :
    tier_fifo_0_io_out_data_count > 14'hd; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_62 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'he :
    tier_fifo_0_io_out_data_count > 14'he; // @[BFS.scala 1354:15]
  wire  _io_cacheable_out_bits_tkeep_T_66 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 14'hf :
    tier_fifo_0_io_out_data_count > 14'hf; // @[BFS.scala 1354:15]
  wire [7:0] io_cacheable_out_bits_tkeep_lo = {_io_cacheable_out_bits_tkeep_T_34,_io_cacheable_out_bits_tkeep_T_30,
    _io_cacheable_out_bits_tkeep_T_26,_io_cacheable_out_bits_tkeep_T_22,_io_cacheable_out_bits_tkeep_T_18,
    _io_cacheable_out_bits_tkeep_T_14,_io_cacheable_out_bits_tkeep_T_10,_io_cacheable_out_bits_tkeep_T_6}; // @[BFS.scala 1355:14]
  wire [15:0] _io_cacheable_out_bits_tkeep_T_67 = {_io_cacheable_out_bits_tkeep_T_66,_io_cacheable_out_bits_tkeep_T_62,
    _io_cacheable_out_bits_tkeep_T_58,_io_cacheable_out_bits_tkeep_T_54,_io_cacheable_out_bits_tkeep_T_50,
    _io_cacheable_out_bits_tkeep_T_46,_io_cacheable_out_bits_tkeep_T_42,_io_cacheable_out_bits_tkeep_T_38,
    io_cacheable_out_bits_tkeep_lo}; // @[BFS.scala 1355:14]
  wire [7:0] _wcount_T_1 = wcount - 8'h1; // @[BFS.scala 1362:22]
  multi_channel_fifo tier_fifo_0 ( // @[BFS.scala 1187:46]
    .clock(tier_fifo_0_clock),
    .reset(tier_fifo_0_reset),
    .io_in_ready(tier_fifo_0_io_in_ready),
    .io_in_valid(tier_fifo_0_io_in_valid),
    .io_in_bits_0_tdata(tier_fifo_0_io_in_bits_0_tdata),
    .io_in_bits_0_tkeep(tier_fifo_0_io_in_bits_0_tkeep),
    .io_in_bits_1_tdata(tier_fifo_0_io_in_bits_1_tdata),
    .io_in_bits_1_tkeep(tier_fifo_0_io_in_bits_1_tkeep),
    .io_in_bits_2_tdata(tier_fifo_0_io_in_bits_2_tdata),
    .io_in_bits_2_tkeep(tier_fifo_0_io_in_bits_2_tkeep),
    .io_in_bits_3_tdata(tier_fifo_0_io_in_bits_3_tdata),
    .io_in_bits_3_tkeep(tier_fifo_0_io_in_bits_3_tkeep),
    .io_in_bits_4_tdata(tier_fifo_0_io_in_bits_4_tdata),
    .io_in_bits_4_tkeep(tier_fifo_0_io_in_bits_4_tkeep),
    .io_in_bits_5_tdata(tier_fifo_0_io_in_bits_5_tdata),
    .io_in_bits_5_tkeep(tier_fifo_0_io_in_bits_5_tkeep),
    .io_in_bits_6_tdata(tier_fifo_0_io_in_bits_6_tdata),
    .io_in_bits_6_tkeep(tier_fifo_0_io_in_bits_6_tkeep),
    .io_in_bits_7_tdata(tier_fifo_0_io_in_bits_7_tdata),
    .io_in_bits_7_tkeep(tier_fifo_0_io_in_bits_7_tkeep),
    .io_in_bits_8_tdata(tier_fifo_0_io_in_bits_8_tdata),
    .io_in_bits_8_tkeep(tier_fifo_0_io_in_bits_8_tkeep),
    .io_in_bits_9_tdata(tier_fifo_0_io_in_bits_9_tdata),
    .io_in_bits_9_tkeep(tier_fifo_0_io_in_bits_9_tkeep),
    .io_in_bits_10_tdata(tier_fifo_0_io_in_bits_10_tdata),
    .io_in_bits_10_tkeep(tier_fifo_0_io_in_bits_10_tkeep),
    .io_in_bits_11_tdata(tier_fifo_0_io_in_bits_11_tdata),
    .io_in_bits_11_tkeep(tier_fifo_0_io_in_bits_11_tkeep),
    .io_in_bits_12_tdata(tier_fifo_0_io_in_bits_12_tdata),
    .io_in_bits_12_tkeep(tier_fifo_0_io_in_bits_12_tkeep),
    .io_in_bits_13_tdata(tier_fifo_0_io_in_bits_13_tdata),
    .io_in_bits_13_tkeep(tier_fifo_0_io_in_bits_13_tkeep),
    .io_in_bits_14_tdata(tier_fifo_0_io_in_bits_14_tdata),
    .io_in_bits_14_tkeep(tier_fifo_0_io_in_bits_14_tkeep),
    .io_in_bits_15_tdata(tier_fifo_0_io_in_bits_15_tdata),
    .io_in_bits_15_tkeep(tier_fifo_0_io_in_bits_15_tkeep),
    .io_out_almost_full(tier_fifo_0_io_out_almost_full),
    .io_out_din(tier_fifo_0_io_out_din),
    .io_out_wr_en(tier_fifo_0_io_out_wr_en),
    .io_out_dout(tier_fifo_0_io_out_dout),
    .io_out_rd_en(tier_fifo_0_io_out_rd_en),
    .io_out_data_count(tier_fifo_0_io_out_data_count),
    .io_out_valid(tier_fifo_0_io_out_valid),
    .io_is_current_tier(tier_fifo_0_io_is_current_tier)
  );
  multi_channel_fifo tier_fifo_1 ( // @[BFS.scala 1187:46]
    .clock(tier_fifo_1_clock),
    .reset(tier_fifo_1_reset),
    .io_in_ready(tier_fifo_1_io_in_ready),
    .io_in_valid(tier_fifo_1_io_in_valid),
    .io_in_bits_0_tdata(tier_fifo_1_io_in_bits_0_tdata),
    .io_in_bits_0_tkeep(tier_fifo_1_io_in_bits_0_tkeep),
    .io_in_bits_1_tdata(tier_fifo_1_io_in_bits_1_tdata),
    .io_in_bits_1_tkeep(tier_fifo_1_io_in_bits_1_tkeep),
    .io_in_bits_2_tdata(tier_fifo_1_io_in_bits_2_tdata),
    .io_in_bits_2_tkeep(tier_fifo_1_io_in_bits_2_tkeep),
    .io_in_bits_3_tdata(tier_fifo_1_io_in_bits_3_tdata),
    .io_in_bits_3_tkeep(tier_fifo_1_io_in_bits_3_tkeep),
    .io_in_bits_4_tdata(tier_fifo_1_io_in_bits_4_tdata),
    .io_in_bits_4_tkeep(tier_fifo_1_io_in_bits_4_tkeep),
    .io_in_bits_5_tdata(tier_fifo_1_io_in_bits_5_tdata),
    .io_in_bits_5_tkeep(tier_fifo_1_io_in_bits_5_tkeep),
    .io_in_bits_6_tdata(tier_fifo_1_io_in_bits_6_tdata),
    .io_in_bits_6_tkeep(tier_fifo_1_io_in_bits_6_tkeep),
    .io_in_bits_7_tdata(tier_fifo_1_io_in_bits_7_tdata),
    .io_in_bits_7_tkeep(tier_fifo_1_io_in_bits_7_tkeep),
    .io_in_bits_8_tdata(tier_fifo_1_io_in_bits_8_tdata),
    .io_in_bits_8_tkeep(tier_fifo_1_io_in_bits_8_tkeep),
    .io_in_bits_9_tdata(tier_fifo_1_io_in_bits_9_tdata),
    .io_in_bits_9_tkeep(tier_fifo_1_io_in_bits_9_tkeep),
    .io_in_bits_10_tdata(tier_fifo_1_io_in_bits_10_tdata),
    .io_in_bits_10_tkeep(tier_fifo_1_io_in_bits_10_tkeep),
    .io_in_bits_11_tdata(tier_fifo_1_io_in_bits_11_tdata),
    .io_in_bits_11_tkeep(tier_fifo_1_io_in_bits_11_tkeep),
    .io_in_bits_12_tdata(tier_fifo_1_io_in_bits_12_tdata),
    .io_in_bits_12_tkeep(tier_fifo_1_io_in_bits_12_tkeep),
    .io_in_bits_13_tdata(tier_fifo_1_io_in_bits_13_tdata),
    .io_in_bits_13_tkeep(tier_fifo_1_io_in_bits_13_tkeep),
    .io_in_bits_14_tdata(tier_fifo_1_io_in_bits_14_tdata),
    .io_in_bits_14_tkeep(tier_fifo_1_io_in_bits_14_tkeep),
    .io_in_bits_15_tdata(tier_fifo_1_io_in_bits_15_tdata),
    .io_in_bits_15_tkeep(tier_fifo_1_io_in_bits_15_tkeep),
    .io_out_almost_full(tier_fifo_1_io_out_almost_full),
    .io_out_din(tier_fifo_1_io_out_din),
    .io_out_wr_en(tier_fifo_1_io_out_wr_en),
    .io_out_dout(tier_fifo_1_io_out_dout),
    .io_out_rd_en(tier_fifo_1_io_out_rd_en),
    .io_out_data_count(tier_fifo_1_io_out_data_count),
    .io_out_valid(tier_fifo_1_io_out_valid),
    .io_is_current_tier(tier_fifo_1_io_is_current_tier)
  );
  multi_channel_fifo_reg_slice in_pipeline_0 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_0_aclk),
    .aresetn(in_pipeline_0_aresetn),
    .s_axis_tdata(in_pipeline_0_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_0_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_0_s_axis_tvalid),
    .s_axis_tready(in_pipeline_0_s_axis_tready),
    .s_axis_tlast(in_pipeline_0_s_axis_tlast),
    .m_axis_tdata(in_pipeline_0_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_0_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_0_m_axis_tvalid),
    .m_axis_tready(in_pipeline_0_m_axis_tready),
    .m_axis_tlast(in_pipeline_0_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_1 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_1_aclk),
    .aresetn(in_pipeline_1_aresetn),
    .s_axis_tdata(in_pipeline_1_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_1_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_1_s_axis_tvalid),
    .s_axis_tready(in_pipeline_1_s_axis_tready),
    .s_axis_tlast(in_pipeline_1_s_axis_tlast),
    .m_axis_tdata(in_pipeline_1_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_1_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_1_m_axis_tvalid),
    .m_axis_tready(in_pipeline_1_m_axis_tready),
    .m_axis_tlast(in_pipeline_1_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_2 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_2_aclk),
    .aresetn(in_pipeline_2_aresetn),
    .s_axis_tdata(in_pipeline_2_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_2_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_2_s_axis_tvalid),
    .s_axis_tready(in_pipeline_2_s_axis_tready),
    .s_axis_tlast(in_pipeline_2_s_axis_tlast),
    .m_axis_tdata(in_pipeline_2_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_2_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_2_m_axis_tvalid),
    .m_axis_tready(in_pipeline_2_m_axis_tready),
    .m_axis_tlast(in_pipeline_2_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_3 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_3_aclk),
    .aresetn(in_pipeline_3_aresetn),
    .s_axis_tdata(in_pipeline_3_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_3_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_3_s_axis_tvalid),
    .s_axis_tready(in_pipeline_3_s_axis_tready),
    .s_axis_tlast(in_pipeline_3_s_axis_tlast),
    .m_axis_tdata(in_pipeline_3_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_3_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_3_m_axis_tvalid),
    .m_axis_tready(in_pipeline_3_m_axis_tready),
    .m_axis_tlast(in_pipeline_3_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_4 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_4_aclk),
    .aresetn(in_pipeline_4_aresetn),
    .s_axis_tdata(in_pipeline_4_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_4_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_4_s_axis_tvalid),
    .s_axis_tready(in_pipeline_4_s_axis_tready),
    .s_axis_tlast(in_pipeline_4_s_axis_tlast),
    .m_axis_tdata(in_pipeline_4_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_4_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_4_m_axis_tvalid),
    .m_axis_tready(in_pipeline_4_m_axis_tready),
    .m_axis_tlast(in_pipeline_4_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_5 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_5_aclk),
    .aresetn(in_pipeline_5_aresetn),
    .s_axis_tdata(in_pipeline_5_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_5_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_5_s_axis_tvalid),
    .s_axis_tready(in_pipeline_5_s_axis_tready),
    .s_axis_tlast(in_pipeline_5_s_axis_tlast),
    .m_axis_tdata(in_pipeline_5_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_5_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_5_m_axis_tvalid),
    .m_axis_tready(in_pipeline_5_m_axis_tready),
    .m_axis_tlast(in_pipeline_5_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_6 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_6_aclk),
    .aresetn(in_pipeline_6_aresetn),
    .s_axis_tdata(in_pipeline_6_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_6_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_6_s_axis_tvalid),
    .s_axis_tready(in_pipeline_6_s_axis_tready),
    .s_axis_tlast(in_pipeline_6_s_axis_tlast),
    .m_axis_tdata(in_pipeline_6_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_6_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_6_m_axis_tvalid),
    .m_axis_tready(in_pipeline_6_m_axis_tready),
    .m_axis_tlast(in_pipeline_6_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_7 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_7_aclk),
    .aresetn(in_pipeline_7_aresetn),
    .s_axis_tdata(in_pipeline_7_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_7_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_7_s_axis_tvalid),
    .s_axis_tready(in_pipeline_7_s_axis_tready),
    .s_axis_tlast(in_pipeline_7_s_axis_tlast),
    .m_axis_tdata(in_pipeline_7_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_7_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_7_m_axis_tvalid),
    .m_axis_tready(in_pipeline_7_m_axis_tready),
    .m_axis_tlast(in_pipeline_7_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_8 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_8_aclk),
    .aresetn(in_pipeline_8_aresetn),
    .s_axis_tdata(in_pipeline_8_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_8_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_8_s_axis_tvalid),
    .s_axis_tready(in_pipeline_8_s_axis_tready),
    .s_axis_tlast(in_pipeline_8_s_axis_tlast),
    .m_axis_tdata(in_pipeline_8_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_8_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_8_m_axis_tvalid),
    .m_axis_tready(in_pipeline_8_m_axis_tready),
    .m_axis_tlast(in_pipeline_8_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_9 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_9_aclk),
    .aresetn(in_pipeline_9_aresetn),
    .s_axis_tdata(in_pipeline_9_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_9_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_9_s_axis_tvalid),
    .s_axis_tready(in_pipeline_9_s_axis_tready),
    .s_axis_tlast(in_pipeline_9_s_axis_tlast),
    .m_axis_tdata(in_pipeline_9_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_9_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_9_m_axis_tvalid),
    .m_axis_tready(in_pipeline_9_m_axis_tready),
    .m_axis_tlast(in_pipeline_9_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_10 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_10_aclk),
    .aresetn(in_pipeline_10_aresetn),
    .s_axis_tdata(in_pipeline_10_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_10_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_10_s_axis_tvalid),
    .s_axis_tready(in_pipeline_10_s_axis_tready),
    .s_axis_tlast(in_pipeline_10_s_axis_tlast),
    .m_axis_tdata(in_pipeline_10_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_10_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_10_m_axis_tvalid),
    .m_axis_tready(in_pipeline_10_m_axis_tready),
    .m_axis_tlast(in_pipeline_10_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_11 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_11_aclk),
    .aresetn(in_pipeline_11_aresetn),
    .s_axis_tdata(in_pipeline_11_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_11_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_11_s_axis_tvalid),
    .s_axis_tready(in_pipeline_11_s_axis_tready),
    .s_axis_tlast(in_pipeline_11_s_axis_tlast),
    .m_axis_tdata(in_pipeline_11_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_11_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_11_m_axis_tvalid),
    .m_axis_tready(in_pipeline_11_m_axis_tready),
    .m_axis_tlast(in_pipeline_11_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_12 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_12_aclk),
    .aresetn(in_pipeline_12_aresetn),
    .s_axis_tdata(in_pipeline_12_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_12_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_12_s_axis_tvalid),
    .s_axis_tready(in_pipeline_12_s_axis_tready),
    .s_axis_tlast(in_pipeline_12_s_axis_tlast),
    .m_axis_tdata(in_pipeline_12_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_12_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_12_m_axis_tvalid),
    .m_axis_tready(in_pipeline_12_m_axis_tready),
    .m_axis_tlast(in_pipeline_12_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_13 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_13_aclk),
    .aresetn(in_pipeline_13_aresetn),
    .s_axis_tdata(in_pipeline_13_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_13_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_13_s_axis_tvalid),
    .s_axis_tready(in_pipeline_13_s_axis_tready),
    .s_axis_tlast(in_pipeline_13_s_axis_tlast),
    .m_axis_tdata(in_pipeline_13_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_13_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_13_m_axis_tvalid),
    .m_axis_tready(in_pipeline_13_m_axis_tready),
    .m_axis_tlast(in_pipeline_13_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_14 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_14_aclk),
    .aresetn(in_pipeline_14_aresetn),
    .s_axis_tdata(in_pipeline_14_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_14_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_14_s_axis_tvalid),
    .s_axis_tready(in_pipeline_14_s_axis_tready),
    .s_axis_tlast(in_pipeline_14_s_axis_tlast),
    .m_axis_tdata(in_pipeline_14_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_14_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_14_m_axis_tvalid),
    .m_axis_tready(in_pipeline_14_m_axis_tready),
    .m_axis_tlast(in_pipeline_14_m_axis_tlast)
  );
  multi_channel_fifo_reg_slice in_pipeline_15 ( // @[BFS.scala 1267:11]
    .aclk(in_pipeline_15_aclk),
    .aresetn(in_pipeline_15_aresetn),
    .s_axis_tdata(in_pipeline_15_s_axis_tdata),
    .s_axis_tkeep(in_pipeline_15_s_axis_tkeep),
    .s_axis_tvalid(in_pipeline_15_s_axis_tvalid),
    .s_axis_tready(in_pipeline_15_s_axis_tready),
    .s_axis_tlast(in_pipeline_15_s_axis_tlast),
    .m_axis_tdata(in_pipeline_15_m_axis_tdata),
    .m_axis_tkeep(in_pipeline_15_m_axis_tkeep),
    .m_axis_tvalid(in_pipeline_15_m_axis_tvalid),
    .m_axis_tready(in_pipeline_15_m_axis_tready),
    .m_axis_tlast(in_pipeline_15_m_axis_tlast)
  );
  assign io_cacheable_out_valid = next_tier_mask[0] ? _io_cacheable_out_valid_T_2 : next_tier_mask[1] &
    _io_cacheable_out_valid_T_5; // @[Mux.scala 98:16]
  assign io_cacheable_out_bits_tdata = _T_5 ? 512'h80000000 : _io_cacheable_out_bits_tdata_T_6; // @[Mux.scala 98:16]
  assign io_cacheable_out_bits_tkeep = _T_5 | _T_14 ? 16'h1 : _io_cacheable_out_bits_tkeep_T_67; // @[BFS.scala 1352:37]
  assign io_cacheable_in_0_ready = in_pipeline_0_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_1_ready = in_pipeline_1_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_2_ready = in_pipeline_2_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_3_ready = in_pipeline_3_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_4_ready = in_pipeline_4_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_5_ready = in_pipeline_5_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_6_ready = in_pipeline_6_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_7_ready = in_pipeline_7_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_8_ready = in_pipeline_8_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_9_ready = in_pipeline_9_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_10_ready = in_pipeline_10_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_11_ready = in_pipeline_11_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_12_ready = in_pipeline_12_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_13_ready = in_pipeline_13_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_14_ready = in_pipeline_14_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_cacheable_in_15_ready = in_pipeline_15_s_axis_tready; // @[BFS.scala 1277:32]
  assign io_ddr_out_0_aw_valid = next_tier_mask[0] ? tier_status_0 == 5'h3 : tier_status_1 == 5'h3; // @[BFS.scala 1370:22]
  assign io_ddr_out_0_aw_bits_awaddr = next_tier_mask[0] ? tier_base_addr_0 : tier_base_addr_1; // @[BFS.scala 1364:28]
  assign io_ddr_out_0_ar_valid = next_tier_mask[0] ? tier_status_1 == 5'h4 : tier_status_0 == 5'h4; // @[BFS.scala 1377:22]
  assign io_ddr_out_0_ar_bits_araddr = next_tier_mask[0] ? tier_base_addr_1 : tier_base_addr_0; // @[BFS.scala 1371:28]
  assign io_ddr_out_0_w_valid = next_tier_mask[0] ? tier_status_0 == 5'h9 : tier_status_1 == 5'h9; // @[BFS.scala 1379:21]
  assign io_ddr_out_0_w_bits_wdata = next_tier_mask[0] ? tier_fifo_0_io_out_dout : tier_fifo_1_io_out_dout; // @[BFS.scala 1378:26]
  assign io_ddr_out_0_w_bits_wlast = wcount == 8'h1; // @[BFS.scala 1380:30]
  assign io_unvisited_size = next_tier_mask[0] ? tier_counter_0 : tier_counter_1; // @[BFS.scala 1343:27]
  assign io_signal_ack = _T_17 | _T_8; // @[BFS.scala 1388:48]
  assign tier_fifo_0_clock = clock;
  assign tier_fifo_0_reset = reset;
  assign tier_fifo_0_io_in_valid = fifo_in_valid_0 | fifo_in_valid_1 | fifo_in_valid_2 | fifo_in_valid_3 |
    fifo_in_valid_4 | fifo_in_valid_5 | fifo_in_valid_6 | fifo_in_valid_7 | fifo_in_valid_8 | fifo_in_valid_9 |
    fifo_in_valid_10 | fifo_in_valid_11 | fifo_in_valid_12 | fifo_in_valid_13 | fifo_in_valid_14 | fifo_in_valid_15; // @[BFS.scala 1313:46]
  assign tier_fifo_0_io_in_bits_0_tdata = _fifo_in_data_T_10 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_190; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_0_tkeep = _fifo_in_data_T_10 ? _steps_T : _fifo_in_valid_T_206; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_1_tdata = _fifo_in_data_T_201 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_381; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_1_tkeep = _fifo_in_data_T_201 ? _steps_T : _fifo_in_valid_T_413; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_2_tdata = _fifo_in_data_T_392 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_572; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_2_tkeep = _fifo_in_data_T_392 ? _steps_T : _fifo_in_valid_T_620; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_3_tdata = _fifo_in_data_T_583 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_763; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_3_tkeep = _fifo_in_data_T_583 ? _steps_T : _fifo_in_valid_T_827; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_4_tdata = _fifo_in_data_T_774 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_954; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_4_tkeep = _fifo_in_data_T_774 ? _steps_T : _fifo_in_valid_T_1034; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_5_tdata = _fifo_in_data_T_965 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1145; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_5_tkeep = _fifo_in_data_T_965 ? _steps_T : _fifo_in_valid_T_1241; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_6_tdata = _fifo_in_data_T_1156 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1336; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_6_tkeep = _fifo_in_data_T_1156 ? _steps_T : _fifo_in_valid_T_1448; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_7_tdata = _fifo_in_data_T_1347 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1527; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_7_tkeep = _fifo_in_data_T_1347 ? _steps_T : _fifo_in_valid_T_1655; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_8_tdata = _fifo_in_data_T_1538 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1718; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_8_tkeep = _fifo_in_data_T_1538 ? _steps_T : _fifo_in_valid_T_1862; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_9_tdata = _fifo_in_data_T_1729 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1909; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_9_tkeep = _fifo_in_data_T_1729 ? _steps_T : _fifo_in_valid_T_2069; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_10_tdata = _fifo_in_data_T_1920 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2100; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_10_tkeep = _fifo_in_data_T_1920 ? _steps_T : _fifo_in_valid_T_2276; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_11_tdata = _fifo_in_data_T_2111 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2291; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_11_tkeep = _fifo_in_data_T_2111 ? _steps_T : _fifo_in_valid_T_2483; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_12_tdata = _fifo_in_data_T_2302 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2482; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_12_tkeep = _fifo_in_data_T_2302 ? _steps_T : _fifo_in_valid_T_2690; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_13_tdata = _fifo_in_data_T_2493 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2673; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_13_tkeep = _fifo_in_data_T_2493 ? _steps_T : _fifo_in_valid_T_2897; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_14_tdata = _fifo_in_data_T_2684 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2864; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_14_tkeep = _fifo_in_data_T_2684 ? _steps_T : _fifo_in_valid_T_3104; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_15_tdata = _fifo_in_data_T_2875 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_3055; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_in_bits_15_tkeep = _fifo_in_data_T_2875 ? _steps_T : _fifo_in_valid_T_3311; // @[Mux.scala 98:16]
  assign tier_fifo_0_io_out_din = next_tier_mask[0] ? 512'h0 : io_ddr_out_0_r_bits_rdata; // @[BFS.scala 1312:26]
  assign tier_fifo_0_io_out_wr_en = next_tier_mask[0] ? 1'h0 : io_ddr_out_0_r_valid; // @[BFS.scala 1311:28]
  assign tier_fifo_0_io_out_rd_en = next_tier_mask[0] ? axi_w_valid & io_ddr_out_0_w_ready :
    _tier_fifo_0_io_out_rd_en_T_4; // @[BFS.scala 1309:28]
  assign tier_fifo_0_io_is_current_tier = ~next_tier_mask[0]; // @[BFS.scala 1321:31]
  assign tier_fifo_1_clock = clock;
  assign tier_fifo_1_reset = reset;
  assign tier_fifo_1_io_in_valid = fifo_in_valid_0 | fifo_in_valid_1 | fifo_in_valid_2 | fifo_in_valid_3 |
    fifo_in_valid_4 | fifo_in_valid_5 | fifo_in_valid_6 | fifo_in_valid_7 | fifo_in_valid_8 | fifo_in_valid_9 |
    fifo_in_valid_10 | fifo_in_valid_11 | fifo_in_valid_12 | fifo_in_valid_13 | fifo_in_valid_14 | fifo_in_valid_15; // @[BFS.scala 1313:46]
  assign tier_fifo_1_io_in_bits_0_tdata = _fifo_in_data_T_10 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_190; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_0_tkeep = _fifo_in_data_T_10 ? _steps_T : _fifo_in_valid_T_206; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_1_tdata = _fifo_in_data_T_201 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_381; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_1_tkeep = _fifo_in_data_T_201 ? _steps_T : _fifo_in_valid_T_413; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_2_tdata = _fifo_in_data_T_392 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_572; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_2_tkeep = _fifo_in_data_T_392 ? _steps_T : _fifo_in_valid_T_620; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_3_tdata = _fifo_in_data_T_583 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_763; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_3_tkeep = _fifo_in_data_T_583 ? _steps_T : _fifo_in_valid_T_827; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_4_tdata = _fifo_in_data_T_774 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_954; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_4_tkeep = _fifo_in_data_T_774 ? _steps_T : _fifo_in_valid_T_1034; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_5_tdata = _fifo_in_data_T_965 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1145; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_5_tkeep = _fifo_in_data_T_965 ? _steps_T : _fifo_in_valid_T_1241; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_6_tdata = _fifo_in_data_T_1156 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1336; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_6_tkeep = _fifo_in_data_T_1156 ? _steps_T : _fifo_in_valid_T_1448; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_7_tdata = _fifo_in_data_T_1347 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1527; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_7_tkeep = _fifo_in_data_T_1347 ? _steps_T : _fifo_in_valid_T_1655; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_8_tdata = _fifo_in_data_T_1538 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1718; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_8_tkeep = _fifo_in_data_T_1538 ? _steps_T : _fifo_in_valid_T_1862; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_9_tdata = _fifo_in_data_T_1729 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_1909; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_9_tkeep = _fifo_in_data_T_1729 ? _steps_T : _fifo_in_valid_T_2069; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_10_tdata = _fifo_in_data_T_1920 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2100; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_10_tkeep = _fifo_in_data_T_1920 ? _steps_T : _fifo_in_valid_T_2276; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_11_tdata = _fifo_in_data_T_2111 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2291; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_11_tkeep = _fifo_in_data_T_2111 ? _steps_T : _fifo_in_valid_T_2483; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_12_tdata = _fifo_in_data_T_2302 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2482; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_12_tkeep = _fifo_in_data_T_2302 ? _steps_T : _fifo_in_valid_T_2690; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_13_tdata = _fifo_in_data_T_2493 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2673; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_13_tkeep = _fifo_in_data_T_2493 ? _steps_T : _fifo_in_valid_T_2897; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_14_tdata = _fifo_in_data_T_2684 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_2864; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_14_tkeep = _fifo_in_data_T_2684 ? _steps_T : _fifo_in_valid_T_3104; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_15_tdata = _fifo_in_data_T_2875 ? in_pipeline_0_m_axis_tdata : _fifo_in_data_T_3055; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_in_bits_15_tkeep = _fifo_in_data_T_2875 ? _steps_T : _fifo_in_valid_T_3311; // @[Mux.scala 98:16]
  assign tier_fifo_1_io_out_din = next_tier_mask[1] ? 512'h0 : io_ddr_out_0_r_bits_rdata; // @[BFS.scala 1312:26]
  assign tier_fifo_1_io_out_wr_en = next_tier_mask[1] ? 1'h0 : io_ddr_out_0_r_valid; // @[BFS.scala 1311:28]
  assign tier_fifo_1_io_out_rd_en = next_tier_mask[1] ? axi_w_valid & io_ddr_out_0_w_ready :
    _tier_fifo_0_io_out_rd_en_T_4; // @[BFS.scala 1309:28]
  assign tier_fifo_1_io_is_current_tier = ~next_tier_mask[1]; // @[BFS.scala 1321:31]
  assign in_pipeline_0_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_0_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_0_s_axis_tdata = io_cacheable_in_0_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_0_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_0_s_axis_tvalid = io_cacheable_in_0_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_0_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_0_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_1_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_1_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_1_s_axis_tdata = io_cacheable_in_1_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_1_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_1_s_axis_tvalid = io_cacheable_in_1_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_1_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_1_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_2_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_2_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_2_s_axis_tdata = io_cacheable_in_2_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_2_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_2_s_axis_tvalid = io_cacheable_in_2_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_2_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_2_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_3_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_3_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_3_s_axis_tdata = io_cacheable_in_3_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_3_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_3_s_axis_tvalid = io_cacheable_in_3_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_3_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_3_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_4_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_4_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_4_s_axis_tdata = io_cacheable_in_4_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_4_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_4_s_axis_tvalid = io_cacheable_in_4_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_4_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_4_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_5_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_5_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_5_s_axis_tdata = io_cacheable_in_5_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_5_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_5_s_axis_tvalid = io_cacheable_in_5_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_5_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_5_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_6_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_6_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_6_s_axis_tdata = io_cacheable_in_6_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_6_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_6_s_axis_tvalid = io_cacheable_in_6_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_6_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_6_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_7_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_7_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_7_s_axis_tdata = io_cacheable_in_7_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_7_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_7_s_axis_tvalid = io_cacheable_in_7_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_7_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_7_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_8_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_8_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_8_s_axis_tdata = io_cacheable_in_8_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_8_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_8_s_axis_tvalid = io_cacheable_in_8_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_8_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_8_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_9_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_9_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_9_s_axis_tdata = io_cacheable_in_9_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_9_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_9_s_axis_tvalid = io_cacheable_in_9_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_9_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_9_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_10_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_10_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_10_s_axis_tdata = io_cacheable_in_10_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_10_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_10_s_axis_tvalid = io_cacheable_in_10_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_10_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_10_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_11_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_11_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_11_s_axis_tdata = io_cacheable_in_11_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_11_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_11_s_axis_tvalid = io_cacheable_in_11_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_11_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_11_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_12_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_12_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_12_s_axis_tdata = io_cacheable_in_12_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_12_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_12_s_axis_tvalid = io_cacheable_in_12_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_12_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_12_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_13_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_13_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_13_s_axis_tdata = io_cacheable_in_13_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_13_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_13_s_axis_tvalid = io_cacheable_in_13_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_13_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_13_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_14_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_14_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_14_s_axis_tdata = io_cacheable_in_14_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_14_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_14_s_axis_tvalid = io_cacheable_in_14_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_14_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_14_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  assign in_pipeline_15_aclk = clock; // @[BFS.scala 1272:32]
  assign in_pipeline_15_aresetn = ~reset; // @[BFS.scala 1273:23]
  assign in_pipeline_15_s_axis_tdata = io_cacheable_in_15_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_pipeline_15_s_axis_tkeep = 4'h1; // @[nf_arm_doce_top.scala 121:11]
  assign in_pipeline_15_s_axis_tvalid = io_cacheable_in_15_valid; // @[BFS.scala 1275:26]
  assign in_pipeline_15_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_pipeline_15_m_axis_tready = next_tier_mask[0] ? tier_fifo_0_io_in_ready : tier_fifo_1_io_in_ready; // @[BFS.scala 1269:24]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1188:29]
      tier_counter_0 <= 32'h0; // @[BFS.scala 1188:29]
    end else if (next_tier_mask[0] & _T_85) begin // @[BFS.scala 1257:97]
      tier_counter_0 <= _tier_counter_0_T_47; // @[BFS.scala 1258:11]
    end else if (_T_35 & io_cacheable_out_ready & io_cacheable_out_valid) begin // @[BFS.scala 1259:89]
      if (tier_fifo_0_io_out_data_count > 14'h10) begin // @[BFS.scala 1260:17]
        tier_counter_0 <= _tier_counter_0_T_50;
      end else begin
        tier_counter_0 <= _tier_counter_0_T_52;
      end
    end
    if (reset) begin // @[BFS.scala 1188:29]
      tier_counter_1 <= 32'h0; // @[BFS.scala 1188:29]
    end else if (next_tier_mask[1] & _T_85) begin // @[BFS.scala 1257:97]
      tier_counter_1 <= _tier_counter_1_T_47; // @[BFS.scala 1258:11]
    end else if (_T_49 & io_cacheable_out_ready & io_cacheable_out_valid) begin // @[BFS.scala 1259:89]
      if (tier_fifo_1_io_out_data_count > 14'h10) begin // @[BFS.scala 1260:17]
        tier_counter_1 <= _tier_counter_1_T_50;
      end else begin
        tier_counter_1 <= _tier_counter_1_T_52;
      end
    end
    if (reset) begin // @[BFS.scala 1206:23]
      status <= 5'h0; // @[BFS.scala 1206:23]
    end else if (io_start & status == 5'h0) begin // @[BFS.scala 1209:40]
      status <= 5'h2; // @[BFS.scala 1210:12]
    end else if (status == 5'h2 & tier_counter_0 == 32'h0) begin // @[BFS.scala 1211:70]
      status <= 5'h5; // @[BFS.scala 1212:12]
    end else if (status == 5'h5 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1213:92]
      status <= 5'h7; // @[BFS.scala 1214:12]
    end else begin
      status <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 1207:28]
      tier_status_0 <= 5'h0; // @[BFS.scala 1207:28]
    end else if (_T_169 & status != 5'h11 & status != 5'h12) begin // @[BFS.scala 1327:69]
      tier_status_0 <= 5'h3; // @[BFS.scala 1328:11]
    end else if (_T_35 & _T_176 & tier_counter_0 != 32'h0 & _T_21) begin // @[BFS.scala 1329:109]
      tier_status_0 <= 5'h4; // @[BFS.scala 1330:11]
    end else if (_axi_aw_valid_T_1 & io_ddr_out_0_aw_ready) begin // @[BFS.scala 1331:53]
      tier_status_0 <= 5'h9; // @[BFS.scala 1332:11]
    end else begin
      tier_status_0 <= _GEN_27;
    end
    if (reset) begin // @[BFS.scala 1207:28]
      tier_status_1 <= 5'h0; // @[BFS.scala 1207:28]
    end else if (_T_199 & status != 5'h11 & status != 5'h12) begin // @[BFS.scala 1327:69]
      tier_status_1 <= 5'h3; // @[BFS.scala 1328:11]
    end else if (_T_49 & _T_206 & tier_counter_1 != 32'h0 & _T_24) begin // @[BFS.scala 1329:109]
      tier_status_1 <= 5'h4; // @[BFS.scala 1330:11]
    end else if (_axi_aw_valid_T_2 & io_ddr_out_0_aw_ready) begin // @[BFS.scala 1331:53]
      tier_status_1 <= 5'h9; // @[BFS.scala 1332:11]
    end else begin
      tier_status_1 <= _GEN_33;
    end
    if (reset) begin // @[BFS.scala 1242:31]
      tier_base_addr_0 <= 64'h0; // @[BFS.scala 1242:31]
    end else if (_T_1 | step_fin) begin // @[BFS.scala 1246:57]
      tier_base_addr_0 <= io_tiers_base_addr_0; // @[BFS.scala 1247:11]
    end else if (next_tier_mask[0] & io_ddr_out_0_aw_ready & axi_aw_valid) begin // @[BFS.scala 1248:86]
      tier_base_addr_0 <= _tier_base_addr_0_T_1; // @[BFS.scala 1249:11]
    end else if (~next_tier_mask[0] & io_ddr_out_0_ar_ready & axi_ar_valid) begin // @[BFS.scala 1250:87]
      tier_base_addr_0 <= _tier_base_addr_0_T_1; // @[BFS.scala 1251:11]
    end
    if (reset) begin // @[BFS.scala 1242:31]
      tier_base_addr_1 <= 64'h0; // @[BFS.scala 1242:31]
    end else if (_T_1 | step_fin) begin // @[BFS.scala 1246:57]
      tier_base_addr_1 <= io_tiers_base_addr_1; // @[BFS.scala 1247:11]
    end else if (next_tier_mask[1] & io_ddr_out_0_aw_ready & axi_aw_valid) begin // @[BFS.scala 1248:86]
      tier_base_addr_1 <= _tier_base_addr_1_T_1; // @[BFS.scala 1249:11]
    end else if (~next_tier_mask[1] & io_ddr_out_0_ar_ready & axi_ar_valid) begin // @[BFS.scala 1250:87]
      tier_base_addr_1 <= _tier_base_addr_1_T_1; // @[BFS.scala 1251:11]
    end
    if (reset) begin // @[BFS.scala 1286:24]
      counter <= 10'h0; // @[BFS.scala 1286:24]
    end else if (steps_15 != 5'h0) begin // @[BFS.scala 1287:39]
      if (_counter_T_1 >= 10'h10) begin // @[BFS.scala 1181:8]
        counter <= _counter_T_6;
      end else begin
        counter <= _counter_T_1;
      end
    end else if (step_fin) begin // @[BFS.scala 1289:88]
      counter <= 10'h0; // @[BFS.scala 1290:13]
    end
    if (reset) begin // @[BFS.scala 1302:30]
      ready_counter <= 32'h0; // @[BFS.scala 1302:30]
    end else if (~fifos_ready & (_steps_T | _steps_T_4 | _steps_T_11 | _steps_T_22 | _steps_T_37 | _steps_T_56 |
      _steps_T_79 | _steps_T_106 | _steps_T_137 | _steps_T_172 | _steps_T_211 | _steps_T_254 | _steps_T_301 |
      _steps_T_352 | _steps_T_407 | _steps_T_466)) begin // @[BFS.scala 1304:97]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 1305:19]
    end
    if (reset) begin // @[BFS.scala 1358:23]
      wcount <= 8'h0; // @[BFS.scala 1358:23]
    end else if (axi_aw_valid & io_ddr_out_0_aw_ready) begin // @[BFS.scala 1359:55]
      wcount <= 8'h10; // @[BFS.scala 1360:12]
    end else if (_tier_fifo_0_io_out_rd_en_T_3) begin // @[BFS.scala 1361:59]
      wcount <= _wcount_T_1; // @[BFS.scala 1362:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tier_counter_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  tier_counter_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  status = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  tier_status_0 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  tier_status_1 = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  tier_base_addr_0 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  tier_base_addr_1 = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  counter = _RAND_7[9:0];
  _RAND_8 = {1{`RANDOM}};
  ready_counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  wcount = _RAND_9[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_arbitrator(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  in_aclk; // @[util.scala 455:18]
  wire  in_aresetn; // @[util.scala 455:18]
  wire [511:0] in_s_axis_tdata; // @[util.scala 455:18]
  wire [63:0] in_s_axis_tkeep; // @[util.scala 455:18]
  wire  in_s_axis_tvalid; // @[util.scala 455:18]
  wire  in_s_axis_tready; // @[util.scala 455:18]
  wire  in_s_axis_tlast; // @[util.scala 455:18]
  wire [511:0] in_m_axis_tdata; // @[util.scala 455:18]
  wire [63:0] in_m_axis_tkeep; // @[util.scala 455:18]
  wire  in_m_axis_tvalid; // @[util.scala 455:18]
  wire  in_m_axis_tready; // @[util.scala 455:18]
  wire  in_m_axis_tlast; // @[util.scala 455:18]
  wire  mid_aclk; // @[util.scala 465:19]
  wire  mid_aresetn; // @[util.scala 465:19]
  wire [511:0] mid_s_axis_tdata; // @[util.scala 465:19]
  wire [63:0] mid_s_axis_tkeep; // @[util.scala 465:19]
  wire  mid_s_axis_tvalid; // @[util.scala 465:19]
  wire  mid_s_axis_tready; // @[util.scala 465:19]
  wire  mid_s_axis_tlast; // @[util.scala 465:19]
  wire [511:0] mid_m_axis_tdata; // @[util.scala 465:19]
  wire [63:0] mid_m_axis_tkeep; // @[util.scala 465:19]
  wire  mid_m_axis_tvalid; // @[util.scala 465:19]
  wire  mid_m_axis_tready; // @[util.scala 465:19]
  wire  mid_m_axis_tlast; // @[util.scala 465:19]
  wire  out_aclk; // @[util.scala 485:19]
  wire  out_aresetn; // @[util.scala 485:19]
  wire [31:0] out_s_axis_tdata; // @[util.scala 485:19]
  wire [3:0] out_s_axis_tkeep; // @[util.scala 485:19]
  wire  out_s_axis_tvalid; // @[util.scala 485:19]
  wire  out_s_axis_tready; // @[util.scala 485:19]
  wire  out_s_axis_tlast; // @[util.scala 485:19]
  wire [31:0] out_m_axis_tdata; // @[util.scala 485:19]
  wire [3:0] out_m_axis_tkeep; // @[util.scala 485:19]
  wire  out_m_axis_tvalid; // @[util.scala 485:19]
  wire  out_m_axis_tready; // @[util.scala 485:19]
  wire  out_m_axis_tlast; // @[util.scala 485:19]
  wire  in_keep_0 = in_m_axis_tkeep[0]; // @[util.scala 463:97]
  wire  in_keep_1 = in_m_axis_tkeep[1]; // @[util.scala 463:97]
  wire  in_keep_2 = in_m_axis_tkeep[2]; // @[util.scala 463:97]
  wire  in_keep_3 = in_m_axis_tkeep[3]; // @[util.scala 463:97]
  wire  in_keep_4 = in_m_axis_tkeep[4]; // @[util.scala 463:97]
  wire  in_keep_5 = in_m_axis_tkeep[5]; // @[util.scala 463:97]
  wire  in_keep_6 = in_m_axis_tkeep[6]; // @[util.scala 463:97]
  wire  in_keep_7 = in_m_axis_tkeep[7]; // @[util.scala 463:97]
  wire  in_keep_8 = in_m_axis_tkeep[8]; // @[util.scala 463:97]
  wire  in_keep_9 = in_m_axis_tkeep[9]; // @[util.scala 463:97]
  wire  in_keep_10 = in_m_axis_tkeep[10]; // @[util.scala 463:97]
  wire  in_keep_11 = in_m_axis_tkeep[11]; // @[util.scala 463:97]
  wire  in_keep_12 = in_m_axis_tkeep[12]; // @[util.scala 463:97]
  wire  in_keep_13 = in_m_axis_tkeep[13]; // @[util.scala 463:97]
  wire  in_keep_14 = in_m_axis_tkeep[14]; // @[util.scala 463:97]
  wire  in_keep_15 = in_m_axis_tkeep[15]; // @[util.scala 463:97]
  wire [4:0] _in_count_WIRE = {{4'd0}, in_keep_0}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_WIRE_1 = {{4'd0}, in_keep_1}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_1 = _in_count_WIRE + _in_count_WIRE_1; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_2 = {{4'd0}, in_keep_2}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_3 = _in_count_T_1 + _in_count_WIRE_2; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_3 = {{4'd0}, in_keep_3}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_5 = _in_count_T_3 + _in_count_WIRE_3; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_4 = {{4'd0}, in_keep_4}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_7 = _in_count_T_5 + _in_count_WIRE_4; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_5 = {{4'd0}, in_keep_5}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_9 = _in_count_T_7 + _in_count_WIRE_5; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_6 = {{4'd0}, in_keep_6}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_11 = _in_count_T_9 + _in_count_WIRE_6; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_7 = {{4'd0}, in_keep_7}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_13 = _in_count_T_11 + _in_count_WIRE_7; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_8 = {{4'd0}, in_keep_8}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_15 = _in_count_T_13 + _in_count_WIRE_8; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_9 = {{4'd0}, in_keep_9}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_17 = _in_count_T_15 + _in_count_WIRE_9; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_10 = {{4'd0}, in_keep_10}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_19 = _in_count_T_17 + _in_count_WIRE_10; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_11 = {{4'd0}, in_keep_11}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_21 = _in_count_T_19 + _in_count_WIRE_11; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_12 = {{4'd0}, in_keep_12}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_23 = _in_count_T_21 + _in_count_WIRE_12; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_13 = {{4'd0}, in_keep_13}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_25 = _in_count_T_23 + _in_count_WIRE_13; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_14 = {{4'd0}, in_keep_14}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_27 = _in_count_T_25 + _in_count_WIRE_14; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_15 = {{4'd0}, in_keep_15}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] in_count = _in_count_T_27 + _in_count_WIRE_15; // @[util.scala 464:82]
  wire [58:0] mid_io_s_axis_tkeep_lo = in_m_axis_tkeep[58:0]; // @[util.scala 472:58]
  wire  keep_0 = mid_m_axis_tkeep[0]; // @[util.scala 476:95]
  wire  keep_1 = mid_m_axis_tkeep[1]; // @[util.scala 476:95]
  wire  keep_2 = mid_m_axis_tkeep[2]; // @[util.scala 476:95]
  wire  keep_3 = mid_m_axis_tkeep[3]; // @[util.scala 476:95]
  wire  keep_4 = mid_m_axis_tkeep[4]; // @[util.scala 476:95]
  wire  keep_5 = mid_m_axis_tkeep[5]; // @[util.scala 476:95]
  wire  keep_6 = mid_m_axis_tkeep[6]; // @[util.scala 476:95]
  wire  keep_7 = mid_m_axis_tkeep[7]; // @[util.scala 476:95]
  wire  keep_8 = mid_m_axis_tkeep[8]; // @[util.scala 476:95]
  wire  keep_9 = mid_m_axis_tkeep[9]; // @[util.scala 476:95]
  wire  keep_10 = mid_m_axis_tkeep[10]; // @[util.scala 476:95]
  wire  keep_11 = mid_m_axis_tkeep[11]; // @[util.scala 476:95]
  wire  keep_12 = mid_m_axis_tkeep[12]; // @[util.scala 476:95]
  wire  keep_13 = mid_m_axis_tkeep[13]; // @[util.scala 476:95]
  wire  keep_14 = mid_m_axis_tkeep[14]; // @[util.scala 476:95]
  wire  keep_15 = mid_m_axis_tkeep[15]; // @[util.scala 476:95]
  reg  index_0; // @[util.scala 477:22]
  reg  index_1; // @[util.scala 477:22]
  reg  index_2; // @[util.scala 477:22]
  reg  index_3; // @[util.scala 477:22]
  reg  index_4; // @[util.scala 477:22]
  reg  index_5; // @[util.scala 477:22]
  reg  index_6; // @[util.scala 477:22]
  reg  index_7; // @[util.scala 477:22]
  reg  index_8; // @[util.scala 477:22]
  reg  index_9; // @[util.scala 477:22]
  reg  index_10; // @[util.scala 477:22]
  reg  index_11; // @[util.scala 477:22]
  reg  index_12; // @[util.scala 477:22]
  reg  index_13; // @[util.scala 477:22]
  reg  index_14; // @[util.scala 477:22]
  reg  index_15; // @[util.scala 477:22]
  wire  ungrant_keep_0 = keep_0 & ~index_0; // @[util.scala 479:22]
  wire  ungrant_keep_1 = keep_1 & ~index_1; // @[util.scala 479:22]
  wire  ungrant_keep_2 = keep_2 & ~index_2; // @[util.scala 479:22]
  wire  ungrant_keep_3 = keep_3 & ~index_3; // @[util.scala 479:22]
  wire  ungrant_keep_4 = keep_4 & ~index_4; // @[util.scala 479:22]
  wire  ungrant_keep_5 = keep_5 & ~index_5; // @[util.scala 479:22]
  wire  ungrant_keep_6 = keep_6 & ~index_6; // @[util.scala 479:22]
  wire  ungrant_keep_7 = keep_7 & ~index_7; // @[util.scala 479:22]
  wire  ungrant_keep_8 = keep_8 & ~index_8; // @[util.scala 479:22]
  wire  ungrant_keep_9 = keep_9 & ~index_9; // @[util.scala 479:22]
  wire  ungrant_keep_10 = keep_10 & ~index_10; // @[util.scala 479:22]
  wire  ungrant_keep_11 = keep_11 & ~index_11; // @[util.scala 479:22]
  wire  ungrant_keep_12 = keep_12 & ~index_12; // @[util.scala 479:22]
  wire  ungrant_keep_13 = keep_13 & ~index_13; // @[util.scala 479:22]
  wire  ungrant_keep_14 = keep_14 & ~index_14; // @[util.scala 479:22]
  wire  ungrant_keep_15 = keep_15 & ~index_15; // @[util.scala 479:22]
  wire  grant_1 = ~ungrant_keep_0; // @[util.scala 363:78]
  wire  grant_2 = ~(ungrant_keep_0 | ungrant_keep_1); // @[util.scala 363:78]
  wire  grant_3 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2); // @[util.scala 363:78]
  wire  grant_4 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3); // @[util.scala 363:78]
  wire  grant_5 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4); // @[util.scala 363:78]
  wire  grant_6 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5)
    ; // @[util.scala 363:78]
  wire  grant_7 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6); // @[util.scala 363:78]
  wire  grant_8 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7); // @[util.scala 363:78]
  wire  grant_9 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8); // @[util.scala 363:78]
  wire  grant_10 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9); // @[util.scala 363:78]
  wire  grant_11 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10); // @[util.scala 363:78]
  wire  grant_12 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10 | ungrant_keep_11); // @[util.scala 363:78]
  wire  grant_13 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10 | ungrant_keep_11 |
    ungrant_keep_12); // @[util.scala 363:78]
  wire  grant_14 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10 | ungrant_keep_11 |
    ungrant_keep_12 | ungrant_keep_13); // @[util.scala 363:78]
  wire  grant_15 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10 | ungrant_keep_11 |
    ungrant_keep_12 | ungrant_keep_13 | ungrant_keep_14); // @[util.scala 363:78]
  wire  choosen_keep_1 = grant_1 & ungrant_keep_1; // @[util.scala 483:22]
  wire  choosen_keep_2 = grant_2 & ungrant_keep_2; // @[util.scala 483:22]
  wire  choosen_keep_3 = grant_3 & ungrant_keep_3; // @[util.scala 483:22]
  wire  choosen_keep_4 = grant_4 & ungrant_keep_4; // @[util.scala 483:22]
  wire  choosen_keep_5 = grant_5 & ungrant_keep_5; // @[util.scala 483:22]
  wire  choosen_keep_6 = grant_6 & ungrant_keep_6; // @[util.scala 483:22]
  wire  choosen_keep_7 = grant_7 & ungrant_keep_7; // @[util.scala 483:22]
  wire  choosen_keep_8 = grant_8 & ungrant_keep_8; // @[util.scala 483:22]
  wire  choosen_keep_9 = grant_9 & ungrant_keep_9; // @[util.scala 483:22]
  wire  choosen_keep_10 = grant_10 & ungrant_keep_10; // @[util.scala 483:22]
  wire  choosen_keep_11 = grant_11 & ungrant_keep_11; // @[util.scala 483:22]
  wire  choosen_keep_12 = grant_12 & ungrant_keep_12; // @[util.scala 483:22]
  wire  choosen_keep_13 = grant_13 & ungrant_keep_13; // @[util.scala 483:22]
  wire  choosen_keep_14 = grant_14 & ungrant_keep_14; // @[util.scala 483:22]
  wire  choosen_keep_15 = grant_15 & ungrant_keep_15; // @[util.scala 483:22]
  wire  _T_1 = mid_m_axis_tvalid; // @[util.scala 491:72]
  wire  _T_4 = out_s_axis_tready; // @[util.scala 493:78]
  wire  _T_5 = out_s_axis_tvalid & out_s_axis_tready; // @[util.scala 493:48]
  reg [4:0] count; // @[util.scala 499:22]
  wire [4:0] next_count = mid_m_axis_tkeep[63:59]; // @[util.scala 500:39]
  wire [4:0] _count_T_1 = next_count - 5'h1; // @[util.scala 503:27]
  wire [4:0] _count_T_3 = count - 5'h1; // @[util.scala 505:22]
  wire [31:0] _out_io_s_axis_tdata_T_16 = ungrant_keep_0 ? mid_m_axis_tdata[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_17 = choosen_keep_1 ? mid_m_axis_tdata[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_18 = choosen_keep_2 ? mid_m_axis_tdata[95:64] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_19 = choosen_keep_3 ? mid_m_axis_tdata[127:96] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_20 = choosen_keep_4 ? mid_m_axis_tdata[159:128] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_21 = choosen_keep_5 ? mid_m_axis_tdata[191:160] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_22 = choosen_keep_6 ? mid_m_axis_tdata[223:192] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_23 = choosen_keep_7 ? mid_m_axis_tdata[255:224] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_24 = choosen_keep_8 ? mid_m_axis_tdata[287:256] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_25 = choosen_keep_9 ? mid_m_axis_tdata[319:288] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_26 = choosen_keep_10 ? mid_m_axis_tdata[351:320] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_27 = choosen_keep_11 ? mid_m_axis_tdata[383:352] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_28 = choosen_keep_12 ? mid_m_axis_tdata[415:384] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_29 = choosen_keep_13 ? mid_m_axis_tdata[447:416] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_30 = choosen_keep_14 ? mid_m_axis_tdata[479:448] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_31 = choosen_keep_15 ? mid_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_32 = _out_io_s_axis_tdata_T_16 | _out_io_s_axis_tdata_T_17; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_33 = _out_io_s_axis_tdata_T_32 | _out_io_s_axis_tdata_T_18; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_34 = _out_io_s_axis_tdata_T_33 | _out_io_s_axis_tdata_T_19; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_35 = _out_io_s_axis_tdata_T_34 | _out_io_s_axis_tdata_T_20; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_36 = _out_io_s_axis_tdata_T_35 | _out_io_s_axis_tdata_T_21; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_37 = _out_io_s_axis_tdata_T_36 | _out_io_s_axis_tdata_T_22; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_38 = _out_io_s_axis_tdata_T_37 | _out_io_s_axis_tdata_T_23; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_39 = _out_io_s_axis_tdata_T_38 | _out_io_s_axis_tdata_T_24; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_40 = _out_io_s_axis_tdata_T_39 | _out_io_s_axis_tdata_T_25; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_41 = _out_io_s_axis_tdata_T_40 | _out_io_s_axis_tdata_T_26; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_42 = _out_io_s_axis_tdata_T_41 | _out_io_s_axis_tdata_T_27; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_43 = _out_io_s_axis_tdata_T_42 | _out_io_s_axis_tdata_T_28; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_44 = _out_io_s_axis_tdata_T_43 | _out_io_s_axis_tdata_T_29; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_45 = _out_io_s_axis_tdata_T_44 | _out_io_s_axis_tdata_T_30; // @[Mux.scala 27:72]
  axis_arbitrator_in_reg_slice_64 in ( // @[util.scala 455:18]
    .aclk(in_aclk),
    .aresetn(in_aresetn),
    .s_axis_tdata(in_s_axis_tdata),
    .s_axis_tkeep(in_s_axis_tkeep),
    .s_axis_tvalid(in_s_axis_tvalid),
    .s_axis_tready(in_s_axis_tready),
    .s_axis_tlast(in_s_axis_tlast),
    .m_axis_tdata(in_m_axis_tdata),
    .m_axis_tkeep(in_m_axis_tkeep),
    .m_axis_tvalid(in_m_axis_tvalid),
    .m_axis_tready(in_m_axis_tready),
    .m_axis_tlast(in_m_axis_tlast)
  );
  axis_arbitrator_in_reg_slice_64 mid ( // @[util.scala 465:19]
    .aclk(mid_aclk),
    .aresetn(mid_aresetn),
    .s_axis_tdata(mid_s_axis_tdata),
    .s_axis_tkeep(mid_s_axis_tkeep),
    .s_axis_tvalid(mid_s_axis_tvalid),
    .s_axis_tready(mid_s_axis_tready),
    .s_axis_tlast(mid_s_axis_tlast),
    .m_axis_tdata(mid_m_axis_tdata),
    .m_axis_tkeep(mid_m_axis_tkeep),
    .m_axis_tvalid(mid_m_axis_tvalid),
    .m_axis_tready(mid_m_axis_tready),
    .m_axis_tlast(mid_m_axis_tlast)
  );
  axis_arbitrator_out_reg_slice_4 out ( // @[util.scala 485:19]
    .aclk(out_aclk),
    .aresetn(out_aresetn),
    .s_axis_tdata(out_s_axis_tdata),
    .s_axis_tkeep(out_s_axis_tkeep),
    .s_axis_tvalid(out_s_axis_tvalid),
    .s_axis_tready(out_s_axis_tready),
    .s_axis_tlast(out_s_axis_tlast),
    .m_axis_tdata(out_m_axis_tdata),
    .m_axis_tkeep(out_m_axis_tkeep),
    .m_axis_tvalid(out_m_axis_tvalid),
    .m_axis_tready(out_m_axis_tready),
    .m_axis_tlast(out_m_axis_tlast)
  );
  assign io_xbar_in_ready = in_s_axis_tready; // @[util.scala 461:20]
  assign io_ddr_out_valid = out_m_axis_tvalid; // @[util.scala 516:20]
  assign io_ddr_out_bits_tdata = out_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign in_aclk = clock; // @[util.scala 457:29]
  assign in_aresetn = ~reset; // @[util.scala 458:20]
  assign in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign in_s_axis_tvalid = io_xbar_in_valid; // @[util.scala 460:23]
  assign in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign in_m_axis_tready = mid_s_axis_tready; // @[util.scala 473:23]
  assign mid_aclk = clock; // @[util.scala 467:30]
  assign mid_aresetn = ~reset; // @[util.scala 468:21]
  assign mid_s_axis_tdata = in_m_axis_tdata; // @[util.scala 470:23]
  assign mid_s_axis_tkeep = {in_count,mid_io_s_axis_tkeep_lo}; // @[Cat.scala 30:58]
  assign mid_s_axis_tvalid = in_m_axis_tvalid; // @[util.scala 469:24]
  assign mid_s_axis_tlast = in_m_axis_tlast; // @[util.scala 471:23]
  assign mid_m_axis_tready = _T_4 & (count == 5'h1 | next_count == 5'h1); // @[util.scala 508:57]
  assign out_aclk = clock; // @[util.scala 486:30]
  assign out_aresetn = ~reset; // @[util.scala 487:21]
  assign out_s_axis_tdata = _out_io_s_axis_tdata_T_45 | _out_io_s_axis_tdata_T_31; // @[Mux.scala 27:72]
  assign out_s_axis_tkeep = 4'h1; // @[util.scala 511:23]
  assign out_s_axis_tvalid = (ungrant_keep_0 | choosen_keep_1 | choosen_keep_2 | choosen_keep_3 | choosen_keep_4 |
    choosen_keep_5 | choosen_keep_6 | choosen_keep_7 | choosen_keep_8 | choosen_keep_9 | choosen_keep_10 |
    choosen_keep_11 | choosen_keep_12 | choosen_keep_13 | choosen_keep_14 | choosen_keep_15) & _T_1; // @[util.scala 510:52]
  assign out_s_axis_tlast = 1'h1; // @[util.scala 512:23]
  assign out_m_axis_tready = io_ddr_out_ready; // @[util.scala 517:24]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 477:22]
      index_0 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_0 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_0 <= index_0 | ungrant_keep_0; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_1 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_1 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_1 <= index_1 | choosen_keep_1; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_2 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_2 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_2 <= index_2 | choosen_keep_2; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_3 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_3 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_3 <= index_3 | choosen_keep_3; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_4 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_4 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_4 <= index_4 | choosen_keep_4; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_5 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_5 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_5 <= index_5 | choosen_keep_5; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_6 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_6 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_6 <= index_6 | choosen_keep_6; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_7 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_7 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_7 <= index_7 | choosen_keep_7; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_8 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_8 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_8 <= index_8 | choosen_keep_8; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_9 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_9 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_9 <= index_9 | choosen_keep_9; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_10 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_10 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_10 <= index_10 | choosen_keep_10; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_11 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_11 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_11 <= index_11 | choosen_keep_11; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_12 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_12 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_12 <= index_12 | choosen_keep_12; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_13 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_13 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_13 <= index_13 | choosen_keep_13; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_14 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_14 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_14 <= index_14 | choosen_keep_14; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_15 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_15 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_15 <= index_15 | choosen_keep_15; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 499:22]
      count <= 5'h0; // @[util.scala 499:22]
    end else if (_T_5) begin // @[util.scala 501:71]
      if (count == 5'h0) begin // @[util.scala 502:24]
        count <= _count_T_1; // @[util.scala 503:13]
      end else begin
        count <= _count_T_3; // @[util.scala 505:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  index_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  index_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  index_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  index_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  index_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  index_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  index_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  index_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  index_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  index_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  index_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  index_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  index_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  index_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  index_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  index_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  count = _RAND_16[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h0; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_1(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h1; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_2(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h2; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_3(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h3; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_4(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h4; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_5(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h5; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_6(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h6; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_7(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h7; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_8(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h8; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_9(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'h9; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_10(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'ha; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_11(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'hb; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_12(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'hc; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_13(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'hd; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_14(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'he; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_15(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 996:22]
  wire  bitmap__clka; // @[BFS.scala 996:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 996:22]
  wire  bitmap__ena; // @[BFS.scala 996:22]
  wire  bitmap__wea; // @[BFS.scala 996:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 996:22]
  wire  bitmap__clkb; // @[BFS.scala 996:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 996:22]
  wire  bitmap__enb; // @[BFS.scala 996:22]
  wire  arbi_clock; // @[BFS.scala 997:20]
  wire  arbi_reset; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 997:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 997:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 997:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 997:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 997:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 997:20]
  wire  scatter_in_aclk; // @[BFS.scala 1022:26]
  wire  scatter_in_aresetn; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 1022:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 1022:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 1022:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 1022:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 1038:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 1038:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 1038:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 1038:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 1051:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1051:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 1051:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 1051:31]
  wire  _filtered_keep_0_T_4 = scatter_in_m_axis_tdata[3:0] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_0_T_5 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_1_T_4 = scatter_in_m_axis_tdata[35:32] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_1_T_5 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_2_T_4 = scatter_in_m_axis_tdata[67:64] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_2_T_5 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_3_T_4 = scatter_in_m_axis_tdata[99:96] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_3_T_5 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_4_T_4 = scatter_in_m_axis_tdata[131:128] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_4_T_5 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_5_T_4 = scatter_in_m_axis_tdata[163:160] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_5_T_5 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_6_T_4 = scatter_in_m_axis_tdata[195:192] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_6_T_5 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_7_T_4 = scatter_in_m_axis_tdata[227:224] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_7_T_5 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_8_T_4 = scatter_in_m_axis_tdata[259:256] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_8_T_5 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_9_T_4 = scatter_in_m_axis_tdata[291:288] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_9_T_5 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_10_T_4 = scatter_in_m_axis_tdata[323:320] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_10_T_5 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_11_T_4 = scatter_in_m_axis_tdata[355:352] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_11_T_5 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_12_T_4 = scatter_in_m_axis_tdata[387:384] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_12_T_5 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_13_T_4 = scatter_in_m_axis_tdata[419:416] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_13_T_5 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_14_T_4 = scatter_in_m_axis_tdata[451:448] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_14_T_5 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[BFS.scala 1032:15]
  wire  _filtered_keep_15_T_4 = scatter_in_m_axis_tdata[483:480] == 4'hf; // @[BFS.scala 1003:39]
  wire  _filtered_keep_15_T_5 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[BFS.scala 1033:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[BFS.scala 1032:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 1044:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 1044:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 1057:47]
  reg  bitmap_wait_valid; // @[BFS.scala 1058:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 1058:28]
  wire  _T = ~halt; // @[BFS.scala 1059:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 1064:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 1064:34]
  wire  _bitmap_write_addr_valid_T_1 = bitmap_wait_bits[30:4] > 27'he7fff; // @[BFS.scala 1017:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[6:4]}; // @[BFS.scala 1019:107 BFS.scala 1019:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = bitmap_wait_bits[30:4] > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 1017:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 1011:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_bits[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_bits[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 1011:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1082:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 1081:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 1070:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 1076:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 1076:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 1067:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 1067:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 1074:56]
  wire [23:0] _GEN_6 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 1074:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_6 | _bitmap_write_data_bits_T_4; // @[BFS.scala 1074:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 1071:14 BFS.scala 1074:28 BFS.scala 1070:34]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = arbi_io_ddr_out_bits_tdata[30:4] - 27'he7fff; // @[BFS.scala 1012:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{3'd0}, arbi_io_ddr_out_bits_tdata[30:7]}; // @[BFS.scala 1013:69 BFS.scala 1013:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = arbi_io_ddr_out_bits_tdata[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_valid_T_5 : _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 1011:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 1078:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 1088:25]
  bitmap_0 bitmap_ ( // @[BFS.scala 996:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 997:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 1022:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 1038:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 1051:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 1027:20]
  assign io_ddr_out_valid = vertex_out_fifo_m_axis_tvalid & ~vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1098:56]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[BFS.scala 1101:25]
  assign io_end = vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]; // @[BFS.scala 1104:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 1096:19]
  assign bitmap__clka = clock; // @[BFS.scala 1094:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 1095:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 1092:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 1093:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 1088:19]
  assign bitmap__clkb = clock; // @[BFS.scala 1089:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 1087:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 1048:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 1086:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 1023:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 1024:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 1026:31]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 1045:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 1039:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 1040:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 1041:34]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 1044:57]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 1043:66]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 1042:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 1049:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 1052:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 1053:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 1091:35]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 1090:36]
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 1097:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 1060:23]
    end
    if (reset) begin // @[BFS.scala 1058:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 1058:28]
    end else if (~halt) begin // @[BFS.scala 1059:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 1061:22]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 1066:29]
    end
    if (reset) begin // @[BFS.scala 1064:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 1064:34]
    end else if (_T) begin // @[BFS.scala 1065:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 1068:28]
    end
    if (reset) begin // @[BFS.scala 1070:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 1070:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 1077:35]
    end
    if (reset) begin // @[BFS.scala 1076:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 1076:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 1079:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_6[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_arbitrator_16(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [127:0] io_xbar_in_bits_tdata,
  input  [3:0]   io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  in_aclk; // @[util.scala 455:18]
  wire  in_aresetn; // @[util.scala 455:18]
  wire [127:0] in_s_axis_tdata; // @[util.scala 455:18]
  wire [15:0] in_s_axis_tkeep; // @[util.scala 455:18]
  wire  in_s_axis_tvalid; // @[util.scala 455:18]
  wire  in_s_axis_tready; // @[util.scala 455:18]
  wire  in_s_axis_tlast; // @[util.scala 455:18]
  wire [127:0] in_m_axis_tdata; // @[util.scala 455:18]
  wire [15:0] in_m_axis_tkeep; // @[util.scala 455:18]
  wire  in_m_axis_tvalid; // @[util.scala 455:18]
  wire  in_m_axis_tready; // @[util.scala 455:18]
  wire  in_m_axis_tlast; // @[util.scala 455:18]
  wire  mid_aclk; // @[util.scala 465:19]
  wire  mid_aresetn; // @[util.scala 465:19]
  wire [127:0] mid_s_axis_tdata; // @[util.scala 465:19]
  wire [15:0] mid_s_axis_tkeep; // @[util.scala 465:19]
  wire  mid_s_axis_tvalid; // @[util.scala 465:19]
  wire  mid_s_axis_tready; // @[util.scala 465:19]
  wire  mid_s_axis_tlast; // @[util.scala 465:19]
  wire [127:0] mid_m_axis_tdata; // @[util.scala 465:19]
  wire [15:0] mid_m_axis_tkeep; // @[util.scala 465:19]
  wire  mid_m_axis_tvalid; // @[util.scala 465:19]
  wire  mid_m_axis_tready; // @[util.scala 465:19]
  wire  mid_m_axis_tlast; // @[util.scala 465:19]
  wire  out_aclk; // @[util.scala 485:19]
  wire  out_aresetn; // @[util.scala 485:19]
  wire [31:0] out_s_axis_tdata; // @[util.scala 485:19]
  wire [3:0] out_s_axis_tkeep; // @[util.scala 485:19]
  wire  out_s_axis_tvalid; // @[util.scala 485:19]
  wire  out_s_axis_tready; // @[util.scala 485:19]
  wire  out_s_axis_tlast; // @[util.scala 485:19]
  wire [31:0] out_m_axis_tdata; // @[util.scala 485:19]
  wire [3:0] out_m_axis_tkeep; // @[util.scala 485:19]
  wire  out_m_axis_tvalid; // @[util.scala 485:19]
  wire  out_m_axis_tready; // @[util.scala 485:19]
  wire  out_m_axis_tlast; // @[util.scala 485:19]
  wire  in_keep_0 = in_m_axis_tkeep[0]; // @[util.scala 463:97]
  wire  in_keep_1 = in_m_axis_tkeep[1]; // @[util.scala 463:97]
  wire  in_keep_2 = in_m_axis_tkeep[2]; // @[util.scala 463:97]
  wire  in_keep_3 = in_m_axis_tkeep[3]; // @[util.scala 463:97]
  wire [2:0] _in_count_WIRE = {{2'd0}, in_keep_0}; // @[util.scala 464:43 util.scala 464:43]
  wire [2:0] _in_count_WIRE_1 = {{2'd0}, in_keep_1}; // @[util.scala 464:43 util.scala 464:43]
  wire [2:0] _in_count_T_1 = _in_count_WIRE + _in_count_WIRE_1; // @[util.scala 464:82]
  wire [2:0] _in_count_WIRE_2 = {{2'd0}, in_keep_2}; // @[util.scala 464:43 util.scala 464:43]
  wire [2:0] _in_count_T_3 = _in_count_T_1 + _in_count_WIRE_2; // @[util.scala 464:82]
  wire [2:0] _in_count_WIRE_3 = {{2'd0}, in_keep_3}; // @[util.scala 464:43 util.scala 464:43]
  wire [2:0] in_count = _in_count_T_3 + _in_count_WIRE_3; // @[util.scala 464:82]
  wire [12:0] mid_io_s_axis_tkeep_lo = in_m_axis_tkeep[12:0]; // @[util.scala 472:58]
  wire  keep_0 = mid_m_axis_tkeep[0]; // @[util.scala 476:95]
  wire  keep_1 = mid_m_axis_tkeep[1]; // @[util.scala 476:95]
  wire  keep_2 = mid_m_axis_tkeep[2]; // @[util.scala 476:95]
  wire  keep_3 = mid_m_axis_tkeep[3]; // @[util.scala 476:95]
  reg  index_0; // @[util.scala 477:22]
  reg  index_1; // @[util.scala 477:22]
  reg  index_2; // @[util.scala 477:22]
  reg  index_3; // @[util.scala 477:22]
  wire  ungrant_keep_0 = keep_0 & ~index_0; // @[util.scala 479:22]
  wire  ungrant_keep_1 = keep_1 & ~index_1; // @[util.scala 479:22]
  wire  ungrant_keep_2 = keep_2 & ~index_2; // @[util.scala 479:22]
  wire  ungrant_keep_3 = keep_3 & ~index_3; // @[util.scala 479:22]
  wire  grant_1 = ~ungrant_keep_0; // @[util.scala 363:78]
  wire  grant_2 = ~(ungrant_keep_0 | ungrant_keep_1); // @[util.scala 363:78]
  wire  grant_3 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2); // @[util.scala 363:78]
  wire  choosen_keep_1 = grant_1 & ungrant_keep_1; // @[util.scala 483:22]
  wire  choosen_keep_2 = grant_2 & ungrant_keep_2; // @[util.scala 483:22]
  wire  choosen_keep_3 = grant_3 & ungrant_keep_3; // @[util.scala 483:22]
  wire  _T_1 = mid_m_axis_tvalid; // @[util.scala 491:72]
  wire  _T_4 = out_s_axis_tready; // @[util.scala 493:78]
  wire  _T_5 = out_s_axis_tvalid & out_s_axis_tready; // @[util.scala 493:48]
  reg [2:0] count; // @[util.scala 499:22]
  wire [2:0] next_count = mid_m_axis_tkeep[15:13]; // @[util.scala 500:39]
  wire [2:0] _count_T_1 = next_count - 3'h1; // @[util.scala 503:27]
  wire [2:0] _count_T_3 = count - 3'h1; // @[util.scala 505:22]
  wire [31:0] _out_io_s_axis_tdata_T_4 = ungrant_keep_0 ? mid_m_axis_tdata[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_5 = choosen_keep_1 ? mid_m_axis_tdata[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_6 = choosen_keep_2 ? mid_m_axis_tdata[95:64] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_7 = choosen_keep_3 ? mid_m_axis_tdata[127:96] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_8 = _out_io_s_axis_tdata_T_4 | _out_io_s_axis_tdata_T_5; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_9 = _out_io_s_axis_tdata_T_8 | _out_io_s_axis_tdata_T_6; // @[Mux.scala 27:72]
  axis_arbitrator_in_reg_slice_16 in ( // @[util.scala 455:18]
    .aclk(in_aclk),
    .aresetn(in_aresetn),
    .s_axis_tdata(in_s_axis_tdata),
    .s_axis_tkeep(in_s_axis_tkeep),
    .s_axis_tvalid(in_s_axis_tvalid),
    .s_axis_tready(in_s_axis_tready),
    .s_axis_tlast(in_s_axis_tlast),
    .m_axis_tdata(in_m_axis_tdata),
    .m_axis_tkeep(in_m_axis_tkeep),
    .m_axis_tvalid(in_m_axis_tvalid),
    .m_axis_tready(in_m_axis_tready),
    .m_axis_tlast(in_m_axis_tlast)
  );
  axis_arbitrator_in_reg_slice_16 mid ( // @[util.scala 465:19]
    .aclk(mid_aclk),
    .aresetn(mid_aresetn),
    .s_axis_tdata(mid_s_axis_tdata),
    .s_axis_tkeep(mid_s_axis_tkeep),
    .s_axis_tvalid(mid_s_axis_tvalid),
    .s_axis_tready(mid_s_axis_tready),
    .s_axis_tlast(mid_s_axis_tlast),
    .m_axis_tdata(mid_m_axis_tdata),
    .m_axis_tkeep(mid_m_axis_tkeep),
    .m_axis_tvalid(mid_m_axis_tvalid),
    .m_axis_tready(mid_m_axis_tready),
    .m_axis_tlast(mid_m_axis_tlast)
  );
  axis_arbitrator_out_reg_slice_4 out ( // @[util.scala 485:19]
    .aclk(out_aclk),
    .aresetn(out_aresetn),
    .s_axis_tdata(out_s_axis_tdata),
    .s_axis_tkeep(out_s_axis_tkeep),
    .s_axis_tvalid(out_s_axis_tvalid),
    .s_axis_tready(out_s_axis_tready),
    .s_axis_tlast(out_s_axis_tlast),
    .m_axis_tdata(out_m_axis_tdata),
    .m_axis_tkeep(out_m_axis_tkeep),
    .m_axis_tvalid(out_m_axis_tvalid),
    .m_axis_tready(out_m_axis_tready),
    .m_axis_tlast(out_m_axis_tlast)
  );
  assign io_xbar_in_ready = in_s_axis_tready; // @[util.scala 461:20]
  assign io_ddr_out_valid = out_m_axis_tvalid; // @[util.scala 516:20]
  assign io_ddr_out_bits_tdata = out_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign in_aclk = clock; // @[util.scala 457:29]
  assign in_aresetn = ~reset; // @[util.scala 458:20]
  assign in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_s_axis_tkeep = {{12'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign in_s_axis_tvalid = io_xbar_in_valid; // @[util.scala 460:23]
  assign in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign in_m_axis_tready = mid_s_axis_tready; // @[util.scala 473:23]
  assign mid_aclk = clock; // @[util.scala 467:30]
  assign mid_aresetn = ~reset; // @[util.scala 468:21]
  assign mid_s_axis_tdata = in_m_axis_tdata; // @[util.scala 470:23]
  assign mid_s_axis_tkeep = {in_count,mid_io_s_axis_tkeep_lo}; // @[Cat.scala 30:58]
  assign mid_s_axis_tvalid = in_m_axis_tvalid; // @[util.scala 469:24]
  assign mid_s_axis_tlast = in_m_axis_tlast; // @[util.scala 471:23]
  assign mid_m_axis_tready = _T_4 & (count == 3'h1 | next_count == 3'h1); // @[util.scala 508:57]
  assign out_aclk = clock; // @[util.scala 486:30]
  assign out_aresetn = ~reset; // @[util.scala 487:21]
  assign out_s_axis_tdata = _out_io_s_axis_tdata_T_9 | _out_io_s_axis_tdata_T_7; // @[Mux.scala 27:72]
  assign out_s_axis_tkeep = 4'h1; // @[util.scala 511:23]
  assign out_s_axis_tvalid = (ungrant_keep_0 | choosen_keep_1 | choosen_keep_2 | choosen_keep_3) & _T_1; // @[util.scala 510:52]
  assign out_s_axis_tlast = 1'h1; // @[util.scala 512:23]
  assign out_m_axis_tready = io_ddr_out_ready; // @[util.scala 517:24]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 477:22]
      index_0 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_0 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_0 <= index_0 | ungrant_keep_0; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_1 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_1 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_1 <= index_1 | choosen_keep_1; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_2 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_2 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_2 <= index_2 | choosen_keep_2; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_3 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_3 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_3 <= index_3 | choosen_keep_3; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 499:22]
      count <= 3'h0; // @[util.scala 499:22]
    end else if (_T_5) begin // @[util.scala 501:71]
      if (count == 3'h0) begin // @[util.scala 502:24]
        count <= _count_T_1; // @[util.scala 503:13]
      end else begin
        count <= _count_T_3; // @[util.scala 505:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  index_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  index_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  index_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  index_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  count = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Gather(
  input          clock,
  input          reset,
  output         io_ddr_in_ready,
  input          io_ddr_in_valid,
  input  [511:0] io_ddr_in_bits_tdata,
  input  [15:0]  io_ddr_in_bits_tkeep,
  input          io_gather_out_0_ready,
  output         io_gather_out_0_valid,
  output [31:0]  io_gather_out_0_bits_tdata,
  input          io_gather_out_1_ready,
  output         io_gather_out_1_valid,
  output [31:0]  io_gather_out_1_bits_tdata,
  input          io_gather_out_2_ready,
  output         io_gather_out_2_valid,
  output [31:0]  io_gather_out_2_bits_tdata,
  input          io_gather_out_3_ready,
  output         io_gather_out_3_valid,
  output [31:0]  io_gather_out_3_bits_tdata,
  input          io_level_cache_out_ready,
  output         io_level_cache_out_valid,
  output [511:0] io_level_cache_out_bits_tdata,
  output [15:0]  io_level_cache_out_bits_tkeep,
  output         io_level_cache_out_bits_tlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  broadcaster_aclk; // @[BFS.scala 330:27]
  wire  broadcaster_aresetn; // @[BFS.scala 330:27]
  wire [511:0] broadcaster_s_axis_tdata; // @[BFS.scala 330:27]
  wire [63:0] broadcaster_s_axis_tkeep; // @[BFS.scala 330:27]
  wire  broadcaster_s_axis_tvalid; // @[BFS.scala 330:27]
  wire  broadcaster_s_axis_tready; // @[BFS.scala 330:27]
  wire  broadcaster_s_axis_tlast; // @[BFS.scala 330:27]
  wire  broadcaster_s_axis_tid; // @[BFS.scala 330:27]
  wire [2559:0] broadcaster_m_axis_tdata; // @[BFS.scala 330:27]
  wire [319:0] broadcaster_m_axis_tkeep; // @[BFS.scala 330:27]
  wire [4:0] broadcaster_m_axis_tvalid; // @[BFS.scala 330:27]
  wire [4:0] broadcaster_m_axis_tready; // @[BFS.scala 330:27]
  wire [4:0] broadcaster_m_axis_tlast; // @[BFS.scala 330:27]
  wire [4:0] broadcaster_m_axis_tid; // @[BFS.scala 330:27]
  wire  v2Apply_fifo_aclk; // @[BFS.scala 337:28]
  wire  v2Apply_fifo_aresetn; // @[BFS.scala 337:28]
  wire [511:0] v2Apply_fifo_s_axis_tdata; // @[BFS.scala 337:28]
  wire [63:0] v2Apply_fifo_s_axis_tkeep; // @[BFS.scala 337:28]
  wire  v2Apply_fifo_s_axis_tvalid; // @[BFS.scala 337:28]
  wire  v2Apply_fifo_s_axis_tready; // @[BFS.scala 337:28]
  wire  v2Apply_fifo_s_axis_tlast; // @[BFS.scala 337:28]
  wire [511:0] v2Apply_fifo_m_axis_tdata; // @[BFS.scala 337:28]
  wire [63:0] v2Apply_fifo_m_axis_tkeep; // @[BFS.scala 337:28]
  wire  v2Apply_fifo_m_axis_tvalid; // @[BFS.scala 337:28]
  wire  v2Apply_fifo_m_axis_tready; // @[BFS.scala 337:28]
  wire  v2Apply_fifo_m_axis_tlast; // @[BFS.scala 337:28]
  wire  v2Broadcast_fifo_0_aclk; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_0_aresetn; // @[BFS.scala 346:16]
  wire [127:0] v2Broadcast_fifo_0_s_axis_tdata; // @[BFS.scala 346:16]
  wire [15:0] v2Broadcast_fifo_0_s_axis_tkeep; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_0_s_axis_tvalid; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_0_s_axis_tready; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_0_s_axis_tlast; // @[BFS.scala 346:16]
  wire [127:0] v2Broadcast_fifo_0_m_axis_tdata; // @[BFS.scala 346:16]
  wire [15:0] v2Broadcast_fifo_0_m_axis_tkeep; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_0_m_axis_tvalid; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_0_m_axis_tready; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_0_m_axis_tlast; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_1_aclk; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_1_aresetn; // @[BFS.scala 346:16]
  wire [127:0] v2Broadcast_fifo_1_s_axis_tdata; // @[BFS.scala 346:16]
  wire [15:0] v2Broadcast_fifo_1_s_axis_tkeep; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_1_s_axis_tvalid; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_1_s_axis_tready; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_1_s_axis_tlast; // @[BFS.scala 346:16]
  wire [127:0] v2Broadcast_fifo_1_m_axis_tdata; // @[BFS.scala 346:16]
  wire [15:0] v2Broadcast_fifo_1_m_axis_tkeep; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_1_m_axis_tvalid; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_1_m_axis_tready; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_1_m_axis_tlast; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_2_aclk; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_2_aresetn; // @[BFS.scala 346:16]
  wire [127:0] v2Broadcast_fifo_2_s_axis_tdata; // @[BFS.scala 346:16]
  wire [15:0] v2Broadcast_fifo_2_s_axis_tkeep; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_2_s_axis_tvalid; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_2_s_axis_tready; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_2_s_axis_tlast; // @[BFS.scala 346:16]
  wire [127:0] v2Broadcast_fifo_2_m_axis_tdata; // @[BFS.scala 346:16]
  wire [15:0] v2Broadcast_fifo_2_m_axis_tkeep; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_2_m_axis_tvalid; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_2_m_axis_tready; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_2_m_axis_tlast; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_3_aclk; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_3_aresetn; // @[BFS.scala 346:16]
  wire [127:0] v2Broadcast_fifo_3_s_axis_tdata; // @[BFS.scala 346:16]
  wire [15:0] v2Broadcast_fifo_3_s_axis_tkeep; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_3_s_axis_tvalid; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_3_s_axis_tready; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_3_s_axis_tlast; // @[BFS.scala 346:16]
  wire [127:0] v2Broadcast_fifo_3_m_axis_tdata; // @[BFS.scala 346:16]
  wire [15:0] v2Broadcast_fifo_3_m_axis_tkeep; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_3_m_axis_tvalid; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_3_m_axis_tready; // @[BFS.scala 346:16]
  wire  v2Broadcast_fifo_3_m_axis_tlast; // @[BFS.scala 346:16]
  wire  v2Broadcast_selecter_0_clock; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_0_reset; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_ready; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_valid; // @[BFS.scala 380:16]
  wire [127:0] v2Broadcast_selecter_0_io_xbar_in_bits_tdata; // @[BFS.scala 380:16]
  wire [3:0] v2Broadcast_selecter_0_io_xbar_in_bits_tkeep; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_bits_tlast; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_0_io_ddr_out_ready; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_0_io_ddr_out_valid; // @[BFS.scala 380:16]
  wire [31:0] v2Broadcast_selecter_0_io_ddr_out_bits_tdata; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_1_clock; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_1_reset; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_ready; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_valid; // @[BFS.scala 380:16]
  wire [127:0] v2Broadcast_selecter_1_io_xbar_in_bits_tdata; // @[BFS.scala 380:16]
  wire [3:0] v2Broadcast_selecter_1_io_xbar_in_bits_tkeep; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_bits_tlast; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_1_io_ddr_out_ready; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_1_io_ddr_out_valid; // @[BFS.scala 380:16]
  wire [31:0] v2Broadcast_selecter_1_io_ddr_out_bits_tdata; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_2_clock; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_2_reset; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_ready; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_valid; // @[BFS.scala 380:16]
  wire [127:0] v2Broadcast_selecter_2_io_xbar_in_bits_tdata; // @[BFS.scala 380:16]
  wire [3:0] v2Broadcast_selecter_2_io_xbar_in_bits_tkeep; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_bits_tlast; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_2_io_ddr_out_ready; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_2_io_ddr_out_valid; // @[BFS.scala 380:16]
  wire [31:0] v2Broadcast_selecter_2_io_ddr_out_bits_tdata; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_3_clock; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_3_reset; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_ready; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_valid; // @[BFS.scala 380:16]
  wire [127:0] v2Broadcast_selecter_3_io_xbar_in_bits_tdata; // @[BFS.scala 380:16]
  wire [3:0] v2Broadcast_selecter_3_io_xbar_in_bits_tkeep; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_bits_tlast; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_3_io_ddr_out_ready; // @[BFS.scala 380:16]
  wire  v2Broadcast_selecter_3_io_ddr_out_valid; // @[BFS.scala 380:16]
  wire [31:0] v2Broadcast_selecter_3_io_ddr_out_bits_tdata; // @[BFS.scala 380:16]
    (*dont_touch = "true" *)reg [31:0] ready_counter; // @[BFS.scala 324:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 327:36]
  wire [63:0] v2Broadcast_fifo_0_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[159:128],broadcaster_m_axis_tdata[31:0]}
    ; // @[BFS.scala 355:16]
  wire [63:0] v2Broadcast_fifo_0_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[415:384],broadcaster_m_axis_tdata[287:
    256]}; // @[BFS.scala 355:16]
  wire  _v2Broadcast_fifo_0_io_s_axis_tvalid_T_29 = broadcaster_m_axis_tkeep[0] | broadcaster_m_axis_tkeep[4] |
    broadcaster_m_axis_tkeep[8] | broadcaster_m_axis_tkeep[12]; // @[BFS.scala 365:17]
  wire [3:0] _v2Broadcast_fifo_0_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[12],broadcaster_m_axis_tkeep[8],
    broadcaster_m_axis_tkeep[4],broadcaster_m_axis_tkeep[0]}; // @[BFS.scala 368:16]
  wire [63:0] v2Broadcast_fifo_1_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[703:672],broadcaster_m_axis_tdata[575:
    544]}; // @[BFS.scala 355:16]
  wire [63:0] v2Broadcast_fifo_1_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[959:928],broadcaster_m_axis_tdata[831:
    800]}; // @[BFS.scala 355:16]
  wire  _v2Broadcast_fifo_1_io_s_axis_tvalid_T_30 = broadcaster_m_axis_tkeep[1] | broadcaster_m_axis_tkeep[5] |
    broadcaster_m_axis_tkeep[9] | broadcaster_m_axis_tkeep[13]; // @[BFS.scala 365:17]
  wire [3:0] _v2Broadcast_fifo_1_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[13],broadcaster_m_axis_tkeep[9],
    broadcaster_m_axis_tkeep[5],broadcaster_m_axis_tkeep[1]}; // @[BFS.scala 368:16]
  wire [63:0] v2Broadcast_fifo_2_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[1247:1216],broadcaster_m_axis_tdata[1119
    :1088]}; // @[BFS.scala 355:16]
  wire [63:0] v2Broadcast_fifo_2_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[1503:1472],broadcaster_m_axis_tdata[1375
    :1344]}; // @[BFS.scala 355:16]
  wire  _v2Broadcast_fifo_2_io_s_axis_tvalid_T_31 = broadcaster_m_axis_tkeep[2] | broadcaster_m_axis_tkeep[6] |
    broadcaster_m_axis_tkeep[10] | broadcaster_m_axis_tkeep[14]; // @[BFS.scala 365:17]
  wire [3:0] _v2Broadcast_fifo_2_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[14],broadcaster_m_axis_tkeep[10],
    broadcaster_m_axis_tkeep[6],broadcaster_m_axis_tkeep[2]}; // @[BFS.scala 368:16]
  wire [63:0] v2Broadcast_fifo_3_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[1791:1760],broadcaster_m_axis_tdata[1663
    :1632]}; // @[BFS.scala 355:16]
  wire [63:0] v2Broadcast_fifo_3_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[2047:2016],broadcaster_m_axis_tdata[1919
    :1888]}; // @[BFS.scala 355:16]
  wire  _v2Broadcast_fifo_3_io_s_axis_tvalid_T_32 = broadcaster_m_axis_tkeep[3] | broadcaster_m_axis_tkeep[7] |
    broadcaster_m_axis_tkeep[11] | broadcaster_m_axis_tkeep[15]; // @[BFS.scala 365:17]
  wire [3:0] _v2Broadcast_fifo_3_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[15],broadcaster_m_axis_tkeep[11],
    broadcaster_m_axis_tkeep[7],broadcaster_m_axis_tkeep[3]}; // @[BFS.scala 368:16]
  wire  _broadcaster_io_m_axis_tready_WIRE_1 = v2Broadcast_fifo_1_s_axis_tready; // @[BFS.scala 373:101 BFS.scala 373:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_0 = v2Broadcast_fifo_0_s_axis_tready; // @[BFS.scala 373:101 BFS.scala 373:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_3 = v2Broadcast_fifo_3_s_axis_tready; // @[BFS.scala 373:101 BFS.scala 373:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_2 = v2Broadcast_fifo_2_s_axis_tready; // @[BFS.scala 373:101 BFS.scala 373:101]
  wire [3:0] broadcaster_io_m_axis_tready_lo_1 = {_broadcaster_io_m_axis_tready_WIRE_3,
    _broadcaster_io_m_axis_tready_WIRE_2,_broadcaster_io_m_axis_tready_WIRE_1,_broadcaster_io_m_axis_tready_WIRE_0}; // @[BFS.scala 373:151]
  wire [63:0] _io_level_cache_out_bits_tkeep_T = v2Apply_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [15:0] _v2Broadcast_selecter_0_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_0_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [15:0] _v2Broadcast_selecter_1_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_1_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [15:0] _v2Broadcast_selecter_2_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_2_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [15:0] _v2Broadcast_selecter_3_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_3_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  gather_broadcaster broadcaster ( // @[BFS.scala 330:27]
    .aclk(broadcaster_aclk),
    .aresetn(broadcaster_aresetn),
    .s_axis_tdata(broadcaster_s_axis_tdata),
    .s_axis_tkeep(broadcaster_s_axis_tkeep),
    .s_axis_tvalid(broadcaster_s_axis_tvalid),
    .s_axis_tready(broadcaster_s_axis_tready),
    .s_axis_tlast(broadcaster_s_axis_tlast),
    .s_axis_tid(broadcaster_s_axis_tid),
    .m_axis_tdata(broadcaster_m_axis_tdata),
    .m_axis_tkeep(broadcaster_m_axis_tkeep),
    .m_axis_tvalid(broadcaster_m_axis_tvalid),
    .m_axis_tready(broadcaster_m_axis_tready),
    .m_axis_tlast(broadcaster_m_axis_tlast),
    .m_axis_tid(broadcaster_m_axis_tid)
  );
  v2A_reg_slice v2Apply_fifo ( // @[BFS.scala 337:28]
    .aclk(v2Apply_fifo_aclk),
    .aresetn(v2Apply_fifo_aresetn),
    .s_axis_tdata(v2Apply_fifo_s_axis_tdata),
    .s_axis_tkeep(v2Apply_fifo_s_axis_tkeep),
    .s_axis_tvalid(v2Apply_fifo_s_axis_tvalid),
    .s_axis_tready(v2Apply_fifo_s_axis_tready),
    .s_axis_tlast(v2Apply_fifo_s_axis_tlast),
    .m_axis_tdata(v2Apply_fifo_m_axis_tdata),
    .m_axis_tkeep(v2Apply_fifo_m_axis_tkeep),
    .m_axis_tvalid(v2Apply_fifo_m_axis_tvalid),
    .m_axis_tready(v2Apply_fifo_m_axis_tready),
    .m_axis_tlast(v2Apply_fifo_m_axis_tlast)
  );
  v2B_reg_slice v2Broadcast_fifo_0 ( // @[BFS.scala 346:16]
    .aclk(v2Broadcast_fifo_0_aclk),
    .aresetn(v2Broadcast_fifo_0_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_0_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_0_s_axis_tkeep),
    .s_axis_tvalid(v2Broadcast_fifo_0_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_0_s_axis_tready),
    .s_axis_tlast(v2Broadcast_fifo_0_s_axis_tlast),
    .m_axis_tdata(v2Broadcast_fifo_0_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_0_m_axis_tkeep),
    .m_axis_tvalid(v2Broadcast_fifo_0_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_0_m_axis_tready),
    .m_axis_tlast(v2Broadcast_fifo_0_m_axis_tlast)
  );
  v2B_reg_slice v2Broadcast_fifo_1 ( // @[BFS.scala 346:16]
    .aclk(v2Broadcast_fifo_1_aclk),
    .aresetn(v2Broadcast_fifo_1_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_1_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_1_s_axis_tkeep),
    .s_axis_tvalid(v2Broadcast_fifo_1_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_1_s_axis_tready),
    .s_axis_tlast(v2Broadcast_fifo_1_s_axis_tlast),
    .m_axis_tdata(v2Broadcast_fifo_1_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_1_m_axis_tkeep),
    .m_axis_tvalid(v2Broadcast_fifo_1_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_1_m_axis_tready),
    .m_axis_tlast(v2Broadcast_fifo_1_m_axis_tlast)
  );
  v2B_reg_slice v2Broadcast_fifo_2 ( // @[BFS.scala 346:16]
    .aclk(v2Broadcast_fifo_2_aclk),
    .aresetn(v2Broadcast_fifo_2_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_2_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_2_s_axis_tkeep),
    .s_axis_tvalid(v2Broadcast_fifo_2_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_2_s_axis_tready),
    .s_axis_tlast(v2Broadcast_fifo_2_s_axis_tlast),
    .m_axis_tdata(v2Broadcast_fifo_2_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_2_m_axis_tkeep),
    .m_axis_tvalid(v2Broadcast_fifo_2_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_2_m_axis_tready),
    .m_axis_tlast(v2Broadcast_fifo_2_m_axis_tlast)
  );
  v2B_reg_slice v2Broadcast_fifo_3 ( // @[BFS.scala 346:16]
    .aclk(v2Broadcast_fifo_3_aclk),
    .aresetn(v2Broadcast_fifo_3_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_3_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_3_s_axis_tkeep),
    .s_axis_tvalid(v2Broadcast_fifo_3_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_3_s_axis_tready),
    .s_axis_tlast(v2Broadcast_fifo_3_s_axis_tlast),
    .m_axis_tdata(v2Broadcast_fifo_3_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_3_m_axis_tkeep),
    .m_axis_tvalid(v2Broadcast_fifo_3_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_3_m_axis_tready),
    .m_axis_tlast(v2Broadcast_fifo_3_m_axis_tlast)
  );
  axis_arbitrator_16 v2Broadcast_selecter_0 ( // @[BFS.scala 380:16]
    .clock(v2Broadcast_selecter_0_clock),
    .reset(v2Broadcast_selecter_0_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_0_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_0_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(v2Broadcast_selecter_0_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(v2Broadcast_selecter_0_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_0_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_0_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_16 v2Broadcast_selecter_1 ( // @[BFS.scala 380:16]
    .clock(v2Broadcast_selecter_1_clock),
    .reset(v2Broadcast_selecter_1_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_1_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_1_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(v2Broadcast_selecter_1_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(v2Broadcast_selecter_1_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_1_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_1_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_16 v2Broadcast_selecter_2 ( // @[BFS.scala 380:16]
    .clock(v2Broadcast_selecter_2_clock),
    .reset(v2Broadcast_selecter_2_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_2_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_2_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(v2Broadcast_selecter_2_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(v2Broadcast_selecter_2_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_2_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_2_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_16 v2Broadcast_selecter_3 ( // @[BFS.scala 380:16]
    .clock(v2Broadcast_selecter_3_clock),
    .reset(v2Broadcast_selecter_3_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_3_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_3_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(v2Broadcast_selecter_3_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(v2Broadcast_selecter_3_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_3_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_3_io_ddr_out_bits_tdata)
  );
  assign io_ddr_in_ready = broadcaster_s_axis_tready; // @[BFS.scala 333:19]
  assign io_gather_out_0_valid = v2Broadcast_selecter_0_io_ddr_out_valid; // @[BFS.scala 387:20]
  assign io_gather_out_0_bits_tdata = v2Broadcast_selecter_0_io_ddr_out_bits_tdata; // @[BFS.scala 387:20]
  assign io_gather_out_1_valid = v2Broadcast_selecter_1_io_ddr_out_valid; // @[BFS.scala 387:20]
  assign io_gather_out_1_bits_tdata = v2Broadcast_selecter_1_io_ddr_out_bits_tdata; // @[BFS.scala 387:20]
  assign io_gather_out_2_valid = v2Broadcast_selecter_2_io_ddr_out_valid; // @[BFS.scala 387:20]
  assign io_gather_out_2_bits_tdata = v2Broadcast_selecter_2_io_ddr_out_bits_tdata; // @[BFS.scala 387:20]
  assign io_gather_out_3_valid = v2Broadcast_selecter_3_io_ddr_out_valid; // @[BFS.scala 387:20]
  assign io_gather_out_3_bits_tdata = v2Broadcast_selecter_3_io_ddr_out_bits_tdata; // @[BFS.scala 387:20]
  assign io_level_cache_out_valid = v2Apply_fifo_m_axis_tvalid; // @[BFS.scala 375:28]
  assign io_level_cache_out_bits_tdata = v2Apply_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_level_cache_out_bits_tkeep = _io_level_cache_out_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_level_cache_out_bits_tlast = v2Apply_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign broadcaster_aclk = clock; // @[BFS.scala 335:38]
  assign broadcaster_aresetn = ~reset; // @[BFS.scala 334:29]
  assign broadcaster_s_axis_tdata = io_ddr_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign broadcaster_s_axis_tkeep = {{48'd0}, io_ddr_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign broadcaster_s_axis_tvalid = io_ddr_in_valid; // @[BFS.scala 332:32]
  assign broadcaster_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign broadcaster_s_axis_tid = 1'h0;
  assign broadcaster_m_axis_tready = {v2Apply_fifo_s_axis_tready,broadcaster_io_m_axis_tready_lo_1}; // @[Cat.scala 30:58]
  assign v2Apply_fifo_aclk = clock; // @[BFS.scala 338:39]
  assign v2Apply_fifo_aresetn = ~reset; // @[BFS.scala 339:30]
  assign v2Apply_fifo_s_axis_tdata = broadcaster_m_axis_tdata[2559:2048]; // @[BFS.scala 340:62]
  assign v2Apply_fifo_s_axis_tkeep = broadcaster_m_axis_tkeep[319:256]; // @[BFS.scala 342:62]
  assign v2Apply_fifo_s_axis_tvalid = broadcaster_m_axis_tvalid[4]; // @[BFS.scala 341:64]
  assign v2Apply_fifo_s_axis_tlast = broadcaster_m_axis_tlast[4]; // @[BFS.scala 343:62]
  assign v2Apply_fifo_m_axis_tready = io_level_cache_out_ready; // @[BFS.scala 376:33]
  assign v2Broadcast_fifo_0_aclk = clock; // @[BFS.scala 351:32]
  assign v2Broadcast_fifo_0_aresetn = ~reset; // @[BFS.scala 350:23]
  assign v2Broadcast_fifo_0_s_axis_tdata = {v2Broadcast_fifo_0_io_s_axis_tdata_hi,v2Broadcast_fifo_0_io_s_axis_tdata_lo}
    ; // @[BFS.scala 355:16]
  assign v2Broadcast_fifo_0_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_0_io_s_axis_tkeep_T_9}; // @[BFS.scala 368:16]
  assign v2Broadcast_fifo_0_s_axis_tvalid = broadcaster_m_axis_tvalid[0] & _v2Broadcast_fifo_0_io_s_axis_tvalid_T_29; // @[BFS.scala 356:61]
  assign v2Broadcast_fifo_0_s_axis_tlast = broadcaster_m_axis_tlast[0]; // @[BFS.scala 369:55]
  assign v2Broadcast_fifo_0_m_axis_tready = v2Broadcast_selecter_0_io_xbar_in_ready; // @[BFS.scala 386:44]
  assign v2Broadcast_fifo_1_aclk = clock; // @[BFS.scala 351:32]
  assign v2Broadcast_fifo_1_aresetn = ~reset; // @[BFS.scala 350:23]
  assign v2Broadcast_fifo_1_s_axis_tdata = {v2Broadcast_fifo_1_io_s_axis_tdata_hi,v2Broadcast_fifo_1_io_s_axis_tdata_lo}
    ; // @[BFS.scala 355:16]
  assign v2Broadcast_fifo_1_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_1_io_s_axis_tkeep_T_9}; // @[BFS.scala 368:16]
  assign v2Broadcast_fifo_1_s_axis_tvalid = broadcaster_m_axis_tvalid[1] & _v2Broadcast_fifo_1_io_s_axis_tvalid_T_30; // @[BFS.scala 356:61]
  assign v2Broadcast_fifo_1_s_axis_tlast = broadcaster_m_axis_tlast[1]; // @[BFS.scala 369:55]
  assign v2Broadcast_fifo_1_m_axis_tready = v2Broadcast_selecter_1_io_xbar_in_ready; // @[BFS.scala 386:44]
  assign v2Broadcast_fifo_2_aclk = clock; // @[BFS.scala 351:32]
  assign v2Broadcast_fifo_2_aresetn = ~reset; // @[BFS.scala 350:23]
  assign v2Broadcast_fifo_2_s_axis_tdata = {v2Broadcast_fifo_2_io_s_axis_tdata_hi,v2Broadcast_fifo_2_io_s_axis_tdata_lo}
    ; // @[BFS.scala 355:16]
  assign v2Broadcast_fifo_2_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_2_io_s_axis_tkeep_T_9}; // @[BFS.scala 368:16]
  assign v2Broadcast_fifo_2_s_axis_tvalid = broadcaster_m_axis_tvalid[2] & _v2Broadcast_fifo_2_io_s_axis_tvalid_T_31; // @[BFS.scala 356:61]
  assign v2Broadcast_fifo_2_s_axis_tlast = broadcaster_m_axis_tlast[2]; // @[BFS.scala 369:55]
  assign v2Broadcast_fifo_2_m_axis_tready = v2Broadcast_selecter_2_io_xbar_in_ready; // @[BFS.scala 386:44]
  assign v2Broadcast_fifo_3_aclk = clock; // @[BFS.scala 351:32]
  assign v2Broadcast_fifo_3_aresetn = ~reset; // @[BFS.scala 350:23]
  assign v2Broadcast_fifo_3_s_axis_tdata = {v2Broadcast_fifo_3_io_s_axis_tdata_hi,v2Broadcast_fifo_3_io_s_axis_tdata_lo}
    ; // @[BFS.scala 355:16]
  assign v2Broadcast_fifo_3_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_3_io_s_axis_tkeep_T_9}; // @[BFS.scala 368:16]
  assign v2Broadcast_fifo_3_s_axis_tvalid = broadcaster_m_axis_tvalid[3] & _v2Broadcast_fifo_3_io_s_axis_tvalid_T_32; // @[BFS.scala 356:61]
  assign v2Broadcast_fifo_3_s_axis_tlast = broadcaster_m_axis_tlast[3]; // @[BFS.scala 369:55]
  assign v2Broadcast_fifo_3_m_axis_tready = v2Broadcast_selecter_3_io_xbar_in_ready; // @[BFS.scala 386:44]
  assign v2Broadcast_selecter_0_clock = clock;
  assign v2Broadcast_selecter_0_reset = reset;
  assign v2Broadcast_selecter_0_io_xbar_in_valid = v2Broadcast_fifo_0_m_axis_tvalid; // @[BFS.scala 384:26]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tdata = v2Broadcast_fifo_0_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_0_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tlast = v2Broadcast_fifo_0_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign v2Broadcast_selecter_0_io_ddr_out_ready = io_gather_out_0_ready; // @[BFS.scala 387:20]
  assign v2Broadcast_selecter_1_clock = clock;
  assign v2Broadcast_selecter_1_reset = reset;
  assign v2Broadcast_selecter_1_io_xbar_in_valid = v2Broadcast_fifo_1_m_axis_tvalid; // @[BFS.scala 384:26]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tdata = v2Broadcast_fifo_1_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_1_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tlast = v2Broadcast_fifo_1_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign v2Broadcast_selecter_1_io_ddr_out_ready = io_gather_out_1_ready; // @[BFS.scala 387:20]
  assign v2Broadcast_selecter_2_clock = clock;
  assign v2Broadcast_selecter_2_reset = reset;
  assign v2Broadcast_selecter_2_io_xbar_in_valid = v2Broadcast_fifo_2_m_axis_tvalid; // @[BFS.scala 384:26]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tdata = v2Broadcast_fifo_2_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_2_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tlast = v2Broadcast_fifo_2_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign v2Broadcast_selecter_2_io_ddr_out_ready = io_gather_out_2_ready; // @[BFS.scala 387:20]
  assign v2Broadcast_selecter_3_clock = clock;
  assign v2Broadcast_selecter_3_reset = reset;
  assign v2Broadcast_selecter_3_io_xbar_in_valid = v2Broadcast_fifo_3_m_axis_tvalid; // @[BFS.scala 384:26]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tdata = v2Broadcast_fifo_3_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_3_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tlast = v2Broadcast_fifo_3_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign v2Broadcast_selecter_3_io_ddr_out_ready = io_gather_out_3_ready; // @[BFS.scala 387:20]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 324:30]
      ready_counter <= 32'h0; // @[BFS.scala 324:30]
    end else if (~io_ddr_in_ready & io_ddr_in_valid) begin // @[BFS.scala 326:66]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 327:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ready_counter = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module URAM_cluster(
  input  [15:0] io_addra,
  input         io_clka,
  input  [47:0] io_dina,
  input         io_wea,
  input  [15:0] io_addrb,
  input         io_clkb,
  output [47:0] io_doutb
);
  wire [11:0] cluster_0_addra; // @[util.scala 123:45]
  wire  cluster_0_clka; // @[util.scala 123:45]
  wire [47:0] cluster_0_dina; // @[util.scala 123:45]
  wire [47:0] cluster_0_douta; // @[util.scala 123:45]
  wire  cluster_0_ena; // @[util.scala 123:45]
  wire  cluster_0_wea; // @[util.scala 123:45]
  wire [11:0] cluster_0_addrb; // @[util.scala 123:45]
  wire  cluster_0_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_0_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_0_doutb; // @[util.scala 123:45]
  wire  cluster_0_enb; // @[util.scala 123:45]
  wire  cluster_0_web; // @[util.scala 123:45]
  wire [11:0] cluster_1_addra; // @[util.scala 123:45]
  wire  cluster_1_clka; // @[util.scala 123:45]
  wire [47:0] cluster_1_dina; // @[util.scala 123:45]
  wire [47:0] cluster_1_douta; // @[util.scala 123:45]
  wire  cluster_1_ena; // @[util.scala 123:45]
  wire  cluster_1_wea; // @[util.scala 123:45]
  wire [11:0] cluster_1_addrb; // @[util.scala 123:45]
  wire  cluster_1_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_1_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_1_doutb; // @[util.scala 123:45]
  wire  cluster_1_enb; // @[util.scala 123:45]
  wire  cluster_1_web; // @[util.scala 123:45]
  wire [11:0] cluster_2_addra; // @[util.scala 123:45]
  wire  cluster_2_clka; // @[util.scala 123:45]
  wire [47:0] cluster_2_dina; // @[util.scala 123:45]
  wire [47:0] cluster_2_douta; // @[util.scala 123:45]
  wire  cluster_2_ena; // @[util.scala 123:45]
  wire  cluster_2_wea; // @[util.scala 123:45]
  wire [11:0] cluster_2_addrb; // @[util.scala 123:45]
  wire  cluster_2_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_2_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_2_doutb; // @[util.scala 123:45]
  wire  cluster_2_enb; // @[util.scala 123:45]
  wire  cluster_2_web; // @[util.scala 123:45]
  wire [11:0] cluster_3_addra; // @[util.scala 123:45]
  wire  cluster_3_clka; // @[util.scala 123:45]
  wire [47:0] cluster_3_dina; // @[util.scala 123:45]
  wire [47:0] cluster_3_douta; // @[util.scala 123:45]
  wire  cluster_3_ena; // @[util.scala 123:45]
  wire  cluster_3_wea; // @[util.scala 123:45]
  wire [11:0] cluster_3_addrb; // @[util.scala 123:45]
  wire  cluster_3_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_3_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_3_doutb; // @[util.scala 123:45]
  wire  cluster_3_enb; // @[util.scala 123:45]
  wire  cluster_3_web; // @[util.scala 123:45]
  wire [11:0] cluster_4_addra; // @[util.scala 123:45]
  wire  cluster_4_clka; // @[util.scala 123:45]
  wire [47:0] cluster_4_dina; // @[util.scala 123:45]
  wire [47:0] cluster_4_douta; // @[util.scala 123:45]
  wire  cluster_4_ena; // @[util.scala 123:45]
  wire  cluster_4_wea; // @[util.scala 123:45]
  wire [11:0] cluster_4_addrb; // @[util.scala 123:45]
  wire  cluster_4_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_4_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_4_doutb; // @[util.scala 123:45]
  wire  cluster_4_enb; // @[util.scala 123:45]
  wire  cluster_4_web; // @[util.scala 123:45]
  wire [11:0] cluster_5_addra; // @[util.scala 123:45]
  wire  cluster_5_clka; // @[util.scala 123:45]
  wire [47:0] cluster_5_dina; // @[util.scala 123:45]
  wire [47:0] cluster_5_douta; // @[util.scala 123:45]
  wire  cluster_5_ena; // @[util.scala 123:45]
  wire  cluster_5_wea; // @[util.scala 123:45]
  wire [11:0] cluster_5_addrb; // @[util.scala 123:45]
  wire  cluster_5_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_5_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_5_doutb; // @[util.scala 123:45]
  wire  cluster_5_enb; // @[util.scala 123:45]
  wire  cluster_5_web; // @[util.scala 123:45]
  wire [11:0] cluster_6_addra; // @[util.scala 123:45]
  wire  cluster_6_clka; // @[util.scala 123:45]
  wire [47:0] cluster_6_dina; // @[util.scala 123:45]
  wire [47:0] cluster_6_douta; // @[util.scala 123:45]
  wire  cluster_6_ena; // @[util.scala 123:45]
  wire  cluster_6_wea; // @[util.scala 123:45]
  wire [11:0] cluster_6_addrb; // @[util.scala 123:45]
  wire  cluster_6_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_6_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_6_doutb; // @[util.scala 123:45]
  wire  cluster_6_enb; // @[util.scala 123:45]
  wire  cluster_6_web; // @[util.scala 123:45]
  wire [11:0] cluster_7_addra; // @[util.scala 123:45]
  wire  cluster_7_clka; // @[util.scala 123:45]
  wire [47:0] cluster_7_dina; // @[util.scala 123:45]
  wire [47:0] cluster_7_douta; // @[util.scala 123:45]
  wire  cluster_7_ena; // @[util.scala 123:45]
  wire  cluster_7_wea; // @[util.scala 123:45]
  wire [11:0] cluster_7_addrb; // @[util.scala 123:45]
  wire  cluster_7_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_7_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_7_doutb; // @[util.scala 123:45]
  wire  cluster_7_enb; // @[util.scala 123:45]
  wire  cluster_7_web; // @[util.scala 123:45]
  wire [11:0] cluster_8_addra; // @[util.scala 123:45]
  wire  cluster_8_clka; // @[util.scala 123:45]
  wire [47:0] cluster_8_dina; // @[util.scala 123:45]
  wire [47:0] cluster_8_douta; // @[util.scala 123:45]
  wire  cluster_8_ena; // @[util.scala 123:45]
  wire  cluster_8_wea; // @[util.scala 123:45]
  wire [11:0] cluster_8_addrb; // @[util.scala 123:45]
  wire  cluster_8_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_8_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_8_doutb; // @[util.scala 123:45]
  wire  cluster_8_enb; // @[util.scala 123:45]
  wire  cluster_8_web; // @[util.scala 123:45]
  wire [11:0] cluster_9_addra; // @[util.scala 123:45]
  wire  cluster_9_clka; // @[util.scala 123:45]
  wire [47:0] cluster_9_dina; // @[util.scala 123:45]
  wire [47:0] cluster_9_douta; // @[util.scala 123:45]
  wire  cluster_9_ena; // @[util.scala 123:45]
  wire  cluster_9_wea; // @[util.scala 123:45]
  wire [11:0] cluster_9_addrb; // @[util.scala 123:45]
  wire  cluster_9_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_9_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_9_doutb; // @[util.scala 123:45]
  wire  cluster_9_enb; // @[util.scala 123:45]
  wire  cluster_9_web; // @[util.scala 123:45]
  wire [11:0] cluster_10_addra; // @[util.scala 123:45]
  wire  cluster_10_clka; // @[util.scala 123:45]
  wire [47:0] cluster_10_dina; // @[util.scala 123:45]
  wire [47:0] cluster_10_douta; // @[util.scala 123:45]
  wire  cluster_10_ena; // @[util.scala 123:45]
  wire  cluster_10_wea; // @[util.scala 123:45]
  wire [11:0] cluster_10_addrb; // @[util.scala 123:45]
  wire  cluster_10_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_10_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_10_doutb; // @[util.scala 123:45]
  wire  cluster_10_enb; // @[util.scala 123:45]
  wire  cluster_10_web; // @[util.scala 123:45]
  wire [11:0] cluster_11_addra; // @[util.scala 123:45]
  wire  cluster_11_clka; // @[util.scala 123:45]
  wire [47:0] cluster_11_dina; // @[util.scala 123:45]
  wire [47:0] cluster_11_douta; // @[util.scala 123:45]
  wire  cluster_11_ena; // @[util.scala 123:45]
  wire  cluster_11_wea; // @[util.scala 123:45]
  wire [11:0] cluster_11_addrb; // @[util.scala 123:45]
  wire  cluster_11_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_11_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_11_doutb; // @[util.scala 123:45]
  wire  cluster_11_enb; // @[util.scala 123:45]
  wire  cluster_11_web; // @[util.scala 123:45]
  wire [11:0] cluster_12_addra; // @[util.scala 123:45]
  wire  cluster_12_clka; // @[util.scala 123:45]
  wire [47:0] cluster_12_dina; // @[util.scala 123:45]
  wire [47:0] cluster_12_douta; // @[util.scala 123:45]
  wire  cluster_12_ena; // @[util.scala 123:45]
  wire  cluster_12_wea; // @[util.scala 123:45]
  wire [11:0] cluster_12_addrb; // @[util.scala 123:45]
  wire  cluster_12_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_12_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_12_doutb; // @[util.scala 123:45]
  wire  cluster_12_enb; // @[util.scala 123:45]
  wire  cluster_12_web; // @[util.scala 123:45]
  wire [11:0] cluster_13_addra; // @[util.scala 123:45]
  wire  cluster_13_clka; // @[util.scala 123:45]
  wire [47:0] cluster_13_dina; // @[util.scala 123:45]
  wire [47:0] cluster_13_douta; // @[util.scala 123:45]
  wire  cluster_13_ena; // @[util.scala 123:45]
  wire  cluster_13_wea; // @[util.scala 123:45]
  wire [11:0] cluster_13_addrb; // @[util.scala 123:45]
  wire  cluster_13_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_13_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_13_doutb; // @[util.scala 123:45]
  wire  cluster_13_enb; // @[util.scala 123:45]
  wire  cluster_13_web; // @[util.scala 123:45]
  wire [11:0] cluster_14_addra; // @[util.scala 123:45]
  wire  cluster_14_clka; // @[util.scala 123:45]
  wire [47:0] cluster_14_dina; // @[util.scala 123:45]
  wire [47:0] cluster_14_douta; // @[util.scala 123:45]
  wire  cluster_14_ena; // @[util.scala 123:45]
  wire  cluster_14_wea; // @[util.scala 123:45]
  wire [11:0] cluster_14_addrb; // @[util.scala 123:45]
  wire  cluster_14_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_14_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_14_doutb; // @[util.scala 123:45]
  wire  cluster_14_enb; // @[util.scala 123:45]
  wire  cluster_14_web; // @[util.scala 123:45]
  wire [11:0] cluster_15_addra; // @[util.scala 123:45]
  wire  cluster_15_clka; // @[util.scala 123:45]
  wire [47:0] cluster_15_dina; // @[util.scala 123:45]
  wire [47:0] cluster_15_douta; // @[util.scala 123:45]
  wire  cluster_15_ena; // @[util.scala 123:45]
  wire  cluster_15_wea; // @[util.scala 123:45]
  wire [11:0] cluster_15_addrb; // @[util.scala 123:45]
  wire  cluster_15_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_15_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_15_doutb; // @[util.scala 123:45]
  wire  cluster_15_enb; // @[util.scala 123:45]
  wire  cluster_15_web; // @[util.scala 123:45]
  wire [15:0] _cluster_0_io_web_T = {{12'd0}, io_addrb[15:12]}; // @[util.scala 137:55]
  wire  _cluster_0_io_web_T_1 = 16'h0 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [15:0] _cluster_0_io_wea_T = {{12'd0}, io_addra[15:12]}; // @[util.scala 138:55]
  wire [47:0] doutb_0 = _cluster_0_io_web_T_1 ? cluster_0_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_1_io_web_T_1 = 16'h1 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_1 = _cluster_1_io_web_T_1 ? cluster_1_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_2_io_web_T_1 = 16'h2 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_2 = _cluster_2_io_web_T_1 ? cluster_2_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_3_io_web_T_1 = 16'h3 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_3 = _cluster_3_io_web_T_1 ? cluster_3_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_4_io_web_T_1 = 16'h4 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_4 = _cluster_4_io_web_T_1 ? cluster_4_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_5_io_web_T_1 = 16'h5 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_5 = _cluster_5_io_web_T_1 ? cluster_5_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_6_io_web_T_1 = 16'h6 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_6 = _cluster_6_io_web_T_1 ? cluster_6_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_7_io_web_T_1 = 16'h7 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_7 = _cluster_7_io_web_T_1 ? cluster_7_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_8_io_web_T_1 = 16'h8 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_8 = _cluster_8_io_web_T_1 ? cluster_8_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_9_io_web_T_1 = 16'h9 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_9 = _cluster_9_io_web_T_1 ? cluster_9_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_10_io_web_T_1 = 16'ha == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_10 = _cluster_10_io_web_T_1 ? cluster_10_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_11_io_web_T_1 = 16'hb == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_11 = _cluster_11_io_web_T_1 ? cluster_11_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_12_io_web_T_1 = 16'hc == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_12 = _cluster_12_io_web_T_1 ? cluster_12_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_13_io_web_T_1 = 16'hd == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_13 = _cluster_13_io_web_T_1 ? cluster_13_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_14_io_web_T_1 = 16'he == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_14 = _cluster_14_io_web_T_1 ? cluster_14_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_15_io_web_T_1 = 16'hf == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_15 = _cluster_15_io_web_T_1 ? cluster_15_doutb : 48'h0; // @[util.scala 139:22]
  wire [47:0] _io_doutb_T = doutb_0 | doutb_1; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_1 = _io_doutb_T | doutb_2; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_2 = _io_doutb_T_1 | doutb_3; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_3 = _io_doutb_T_2 | doutb_4; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_4 = _io_doutb_T_3 | doutb_5; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_5 = _io_doutb_T_4 | doutb_6; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_6 = _io_doutb_T_5 | doutb_7; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_7 = _io_doutb_T_6 | doutb_8; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_8 = _io_doutb_T_7 | doutb_9; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_9 = _io_doutb_T_8 | doutb_10; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_10 = _io_doutb_T_9 | doutb_11; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_11 = _io_doutb_T_10 | doutb_12; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_12 = _io_doutb_T_11 | doutb_13; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_13 = _io_doutb_T_12 | doutb_14; // @[util.scala 144:29]
  URAM cluster_0 ( // @[util.scala 123:45]
    .addra(cluster_0_addra),
    .clka(cluster_0_clka),
    .dina(cluster_0_dina),
    .douta(cluster_0_douta),
    .ena(cluster_0_ena),
    .wea(cluster_0_wea),
    .addrb(cluster_0_addrb),
    .clkb(cluster_0_clkb),
    .dinb(cluster_0_dinb),
    .doutb(cluster_0_doutb),
    .enb(cluster_0_enb),
    .web(cluster_0_web)
  );
  URAM cluster_1 ( // @[util.scala 123:45]
    .addra(cluster_1_addra),
    .clka(cluster_1_clka),
    .dina(cluster_1_dina),
    .douta(cluster_1_douta),
    .ena(cluster_1_ena),
    .wea(cluster_1_wea),
    .addrb(cluster_1_addrb),
    .clkb(cluster_1_clkb),
    .dinb(cluster_1_dinb),
    .doutb(cluster_1_doutb),
    .enb(cluster_1_enb),
    .web(cluster_1_web)
  );
  URAM cluster_2 ( // @[util.scala 123:45]
    .addra(cluster_2_addra),
    .clka(cluster_2_clka),
    .dina(cluster_2_dina),
    .douta(cluster_2_douta),
    .ena(cluster_2_ena),
    .wea(cluster_2_wea),
    .addrb(cluster_2_addrb),
    .clkb(cluster_2_clkb),
    .dinb(cluster_2_dinb),
    .doutb(cluster_2_doutb),
    .enb(cluster_2_enb),
    .web(cluster_2_web)
  );
  URAM cluster_3 ( // @[util.scala 123:45]
    .addra(cluster_3_addra),
    .clka(cluster_3_clka),
    .dina(cluster_3_dina),
    .douta(cluster_3_douta),
    .ena(cluster_3_ena),
    .wea(cluster_3_wea),
    .addrb(cluster_3_addrb),
    .clkb(cluster_3_clkb),
    .dinb(cluster_3_dinb),
    .doutb(cluster_3_doutb),
    .enb(cluster_3_enb),
    .web(cluster_3_web)
  );
  URAM cluster_4 ( // @[util.scala 123:45]
    .addra(cluster_4_addra),
    .clka(cluster_4_clka),
    .dina(cluster_4_dina),
    .douta(cluster_4_douta),
    .ena(cluster_4_ena),
    .wea(cluster_4_wea),
    .addrb(cluster_4_addrb),
    .clkb(cluster_4_clkb),
    .dinb(cluster_4_dinb),
    .doutb(cluster_4_doutb),
    .enb(cluster_4_enb),
    .web(cluster_4_web)
  );
  URAM cluster_5 ( // @[util.scala 123:45]
    .addra(cluster_5_addra),
    .clka(cluster_5_clka),
    .dina(cluster_5_dina),
    .douta(cluster_5_douta),
    .ena(cluster_5_ena),
    .wea(cluster_5_wea),
    .addrb(cluster_5_addrb),
    .clkb(cluster_5_clkb),
    .dinb(cluster_5_dinb),
    .doutb(cluster_5_doutb),
    .enb(cluster_5_enb),
    .web(cluster_5_web)
  );
  URAM cluster_6 ( // @[util.scala 123:45]
    .addra(cluster_6_addra),
    .clka(cluster_6_clka),
    .dina(cluster_6_dina),
    .douta(cluster_6_douta),
    .ena(cluster_6_ena),
    .wea(cluster_6_wea),
    .addrb(cluster_6_addrb),
    .clkb(cluster_6_clkb),
    .dinb(cluster_6_dinb),
    .doutb(cluster_6_doutb),
    .enb(cluster_6_enb),
    .web(cluster_6_web)
  );
  URAM cluster_7 ( // @[util.scala 123:45]
    .addra(cluster_7_addra),
    .clka(cluster_7_clka),
    .dina(cluster_7_dina),
    .douta(cluster_7_douta),
    .ena(cluster_7_ena),
    .wea(cluster_7_wea),
    .addrb(cluster_7_addrb),
    .clkb(cluster_7_clkb),
    .dinb(cluster_7_dinb),
    .doutb(cluster_7_doutb),
    .enb(cluster_7_enb),
    .web(cluster_7_web)
  );
  URAM cluster_8 ( // @[util.scala 123:45]
    .addra(cluster_8_addra),
    .clka(cluster_8_clka),
    .dina(cluster_8_dina),
    .douta(cluster_8_douta),
    .ena(cluster_8_ena),
    .wea(cluster_8_wea),
    .addrb(cluster_8_addrb),
    .clkb(cluster_8_clkb),
    .dinb(cluster_8_dinb),
    .doutb(cluster_8_doutb),
    .enb(cluster_8_enb),
    .web(cluster_8_web)
  );
  URAM cluster_9 ( // @[util.scala 123:45]
    .addra(cluster_9_addra),
    .clka(cluster_9_clka),
    .dina(cluster_9_dina),
    .douta(cluster_9_douta),
    .ena(cluster_9_ena),
    .wea(cluster_9_wea),
    .addrb(cluster_9_addrb),
    .clkb(cluster_9_clkb),
    .dinb(cluster_9_dinb),
    .doutb(cluster_9_doutb),
    .enb(cluster_9_enb),
    .web(cluster_9_web)
  );
  URAM cluster_10 ( // @[util.scala 123:45]
    .addra(cluster_10_addra),
    .clka(cluster_10_clka),
    .dina(cluster_10_dina),
    .douta(cluster_10_douta),
    .ena(cluster_10_ena),
    .wea(cluster_10_wea),
    .addrb(cluster_10_addrb),
    .clkb(cluster_10_clkb),
    .dinb(cluster_10_dinb),
    .doutb(cluster_10_doutb),
    .enb(cluster_10_enb),
    .web(cluster_10_web)
  );
  URAM cluster_11 ( // @[util.scala 123:45]
    .addra(cluster_11_addra),
    .clka(cluster_11_clka),
    .dina(cluster_11_dina),
    .douta(cluster_11_douta),
    .ena(cluster_11_ena),
    .wea(cluster_11_wea),
    .addrb(cluster_11_addrb),
    .clkb(cluster_11_clkb),
    .dinb(cluster_11_dinb),
    .doutb(cluster_11_doutb),
    .enb(cluster_11_enb),
    .web(cluster_11_web)
  );
  URAM cluster_12 ( // @[util.scala 123:45]
    .addra(cluster_12_addra),
    .clka(cluster_12_clka),
    .dina(cluster_12_dina),
    .douta(cluster_12_douta),
    .ena(cluster_12_ena),
    .wea(cluster_12_wea),
    .addrb(cluster_12_addrb),
    .clkb(cluster_12_clkb),
    .dinb(cluster_12_dinb),
    .doutb(cluster_12_doutb),
    .enb(cluster_12_enb),
    .web(cluster_12_web)
  );
  URAM cluster_13 ( // @[util.scala 123:45]
    .addra(cluster_13_addra),
    .clka(cluster_13_clka),
    .dina(cluster_13_dina),
    .douta(cluster_13_douta),
    .ena(cluster_13_ena),
    .wea(cluster_13_wea),
    .addrb(cluster_13_addrb),
    .clkb(cluster_13_clkb),
    .dinb(cluster_13_dinb),
    .doutb(cluster_13_doutb),
    .enb(cluster_13_enb),
    .web(cluster_13_web)
  );
  URAM cluster_14 ( // @[util.scala 123:45]
    .addra(cluster_14_addra),
    .clka(cluster_14_clka),
    .dina(cluster_14_dina),
    .douta(cluster_14_douta),
    .ena(cluster_14_ena),
    .wea(cluster_14_wea),
    .addrb(cluster_14_addrb),
    .clkb(cluster_14_clkb),
    .dinb(cluster_14_dinb),
    .doutb(cluster_14_doutb),
    .enb(cluster_14_enb),
    .web(cluster_14_web)
  );
  URAM cluster_15 ( // @[util.scala 123:45]
    .addra(cluster_15_addra),
    .clka(cluster_15_clka),
    .dina(cluster_15_dina),
    .douta(cluster_15_douta),
    .ena(cluster_15_ena),
    .wea(cluster_15_wea),
    .addrb(cluster_15_addrb),
    .clkb(cluster_15_clkb),
    .dinb(cluster_15_dinb),
    .doutb(cluster_15_doutb),
    .enb(cluster_15_enb),
    .web(cluster_15_web)
  );
  assign io_doutb = _io_doutb_T_13 | doutb_15; // @[util.scala 144:29]
  assign cluster_0_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_0_clka = io_clka; // @[util.scala 130:17]
  assign cluster_0_dina = io_dina; // @[util.scala 134:17]
  assign cluster_0_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_0_wea = io_wea & 16'h0 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_0_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_0_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_0_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_0_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_0_web = 1'h0; // @[util.scala 137:26]
  assign cluster_1_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_1_clka = io_clka; // @[util.scala 130:17]
  assign cluster_1_dina = io_dina; // @[util.scala 134:17]
  assign cluster_1_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_1_wea = io_wea & 16'h1 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_1_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_1_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_1_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_1_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_1_web = 1'h0; // @[util.scala 137:26]
  assign cluster_2_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_2_clka = io_clka; // @[util.scala 130:17]
  assign cluster_2_dina = io_dina; // @[util.scala 134:17]
  assign cluster_2_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_2_wea = io_wea & 16'h2 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_2_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_2_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_2_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_2_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_2_web = 1'h0; // @[util.scala 137:26]
  assign cluster_3_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_3_clka = io_clka; // @[util.scala 130:17]
  assign cluster_3_dina = io_dina; // @[util.scala 134:17]
  assign cluster_3_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_3_wea = io_wea & 16'h3 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_3_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_3_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_3_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_3_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_3_web = 1'h0; // @[util.scala 137:26]
  assign cluster_4_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_4_clka = io_clka; // @[util.scala 130:17]
  assign cluster_4_dina = io_dina; // @[util.scala 134:17]
  assign cluster_4_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_4_wea = io_wea & 16'h4 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_4_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_4_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_4_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_4_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_4_web = 1'h0; // @[util.scala 137:26]
  assign cluster_5_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_5_clka = io_clka; // @[util.scala 130:17]
  assign cluster_5_dina = io_dina; // @[util.scala 134:17]
  assign cluster_5_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_5_wea = io_wea & 16'h5 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_5_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_5_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_5_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_5_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_5_web = 1'h0; // @[util.scala 137:26]
  assign cluster_6_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_6_clka = io_clka; // @[util.scala 130:17]
  assign cluster_6_dina = io_dina; // @[util.scala 134:17]
  assign cluster_6_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_6_wea = io_wea & 16'h6 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_6_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_6_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_6_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_6_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_6_web = 1'h0; // @[util.scala 137:26]
  assign cluster_7_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_7_clka = io_clka; // @[util.scala 130:17]
  assign cluster_7_dina = io_dina; // @[util.scala 134:17]
  assign cluster_7_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_7_wea = io_wea & 16'h7 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_7_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_7_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_7_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_7_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_7_web = 1'h0; // @[util.scala 137:26]
  assign cluster_8_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_8_clka = io_clka; // @[util.scala 130:17]
  assign cluster_8_dina = io_dina; // @[util.scala 134:17]
  assign cluster_8_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_8_wea = io_wea & 16'h8 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_8_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_8_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_8_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_8_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_8_web = 1'h0; // @[util.scala 137:26]
  assign cluster_9_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_9_clka = io_clka; // @[util.scala 130:17]
  assign cluster_9_dina = io_dina; // @[util.scala 134:17]
  assign cluster_9_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_9_wea = io_wea & 16'h9 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_9_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_9_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_9_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_9_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_9_web = 1'h0; // @[util.scala 137:26]
  assign cluster_10_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_10_clka = io_clka; // @[util.scala 130:17]
  assign cluster_10_dina = io_dina; // @[util.scala 134:17]
  assign cluster_10_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_10_wea = io_wea & 16'ha == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_10_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_10_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_10_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_10_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_10_web = 1'h0; // @[util.scala 137:26]
  assign cluster_11_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_11_clka = io_clka; // @[util.scala 130:17]
  assign cluster_11_dina = io_dina; // @[util.scala 134:17]
  assign cluster_11_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_11_wea = io_wea & 16'hb == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_11_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_11_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_11_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_11_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_11_web = 1'h0; // @[util.scala 137:26]
  assign cluster_12_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_12_clka = io_clka; // @[util.scala 130:17]
  assign cluster_12_dina = io_dina; // @[util.scala 134:17]
  assign cluster_12_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_12_wea = io_wea & 16'hc == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_12_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_12_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_12_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_12_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_12_web = 1'h0; // @[util.scala 137:26]
  assign cluster_13_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_13_clka = io_clka; // @[util.scala 130:17]
  assign cluster_13_dina = io_dina; // @[util.scala 134:17]
  assign cluster_13_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_13_wea = io_wea & 16'hd == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_13_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_13_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_13_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_13_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_13_web = 1'h0; // @[util.scala 137:26]
  assign cluster_14_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_14_clka = io_clka; // @[util.scala 130:17]
  assign cluster_14_dina = io_dina; // @[util.scala 134:17]
  assign cluster_14_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_14_wea = io_wea & 16'he == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_14_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_14_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_14_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_14_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_14_web = 1'h0; // @[util.scala 137:26]
  assign cluster_15_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_15_clka = io_clka; // @[util.scala 130:17]
  assign cluster_15_dina = io_dina; // @[util.scala 134:17]
  assign cluster_15_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_15_wea = io_wea & 16'hf == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_15_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_15_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_15_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_15_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_15_web = 1'h0; // @[util.scala 137:26]
endmodule
module WB_engine(
  input          clock,
  input          reset,
  input          io_axi_ddr_aw_ready,
  output         io_axi_ddr_aw_valid,
  output [63:0]  io_axi_ddr_aw_bits_awaddr,
  output [5:0]   io_axi_ddr_aw_bits_awid,
  input          io_axi_ddr_w_ready,
  output         io_axi_ddr_w_valid,
  output [127:0] io_axi_ddr_w_bits_wdata,
  output [15:0]  io_axi_ddr_w_bits_wstrb,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [31:0]  io_xbar_in_bits_tdata,
  input  [63:0]  io_level_base_addr,
  input  [31:0]  io_level,
  output         io_end,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] buffer_io_addra; // @[BFS.scala 25:22]
  wire  buffer_io_clka; // @[BFS.scala 25:22]
  wire [47:0] buffer_io_dina; // @[BFS.scala 25:22]
  wire  buffer_io_wea; // @[BFS.scala 25:22]
  wire [15:0] buffer_io_addrb; // @[BFS.scala 25:22]
  wire  buffer_io_clkb; // @[BFS.scala 25:22]
  wire [47:0] buffer_io_doutb; // @[BFS.scala 25:22]
  wire [9:0] region_counter__addra; // @[BFS.scala 26:30]
  wire  region_counter__clka; // @[BFS.scala 26:30]
  wire [8:0] region_counter__dina; // @[BFS.scala 26:30]
  wire  region_counter__ena; // @[BFS.scala 26:30]
  wire  region_counter__wea; // @[BFS.scala 26:30]
  wire [9:0] region_counter__addrb; // @[BFS.scala 26:30]
  wire  region_counter__clkb; // @[BFS.scala 26:30]
  wire [8:0] region_counter__doutb; // @[BFS.scala 26:30]
  wire  region_counter__enb; // @[BFS.scala 26:30]
  wire  region_counter_doutb_forward_aclk; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_aresetn; // @[BFS.scala 60:44]
  wire [15:0] region_counter_doutb_forward_s_axis_tdata; // @[BFS.scala 60:44]
  wire [1:0] region_counter_doutb_forward_s_axis_tkeep; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tvalid; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tready; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tlast; // @[BFS.scala 60:44]
  wire [15:0] region_counter_doutb_forward_m_axis_tdata; // @[BFS.scala 60:44]
  wire [1:0] region_counter_doutb_forward_m_axis_tkeep; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tvalid; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tready; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tlast; // @[BFS.scala 60:44]
  wire  pipeline_1_aclk; // @[BFS.scala 64:26]
  wire  pipeline_1_aresetn; // @[BFS.scala 64:26]
  wire [31:0] pipeline_1_s_axis_tdata; // @[BFS.scala 64:26]
  wire [3:0] pipeline_1_s_axis_tkeep; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tvalid; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tready; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tlast; // @[BFS.scala 64:26]
  wire [31:0] pipeline_1_m_axis_tdata; // @[BFS.scala 64:26]
  wire [3:0] pipeline_1_m_axis_tkeep; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tvalid; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tready; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tlast; // @[BFS.scala 64:26]
  wire  aw_buffer_full; // @[BFS.scala 102:25]
  wire [63:0] aw_buffer_din; // @[BFS.scala 102:25]
  wire  aw_buffer_wr_en; // @[BFS.scala 102:25]
  wire  aw_buffer_empty; // @[BFS.scala 102:25]
  wire [63:0] aw_buffer_dout; // @[BFS.scala 102:25]
  wire  aw_buffer_rd_en; // @[BFS.scala 102:25]
  wire [5:0] aw_buffer_data_count; // @[BFS.scala 102:25]
  wire  aw_buffer_clk; // @[BFS.scala 102:25]
  wire  aw_buffer_srst; // @[BFS.scala 102:25]
  wire  aw_buffer_valid; // @[BFS.scala 102:25]
  wire  w_buffer_full; // @[BFS.scala 103:24]
  wire [63:0] w_buffer_din; // @[BFS.scala 103:24]
  wire  w_buffer_wr_en; // @[BFS.scala 103:24]
  wire  w_buffer_empty; // @[BFS.scala 103:24]
  wire [63:0] w_buffer_dout; // @[BFS.scala 103:24]
  wire  w_buffer_rd_en; // @[BFS.scala 103:24]
  wire [5:0] w_buffer_data_count; // @[BFS.scala 103:24]
  wire  w_buffer_clk; // @[BFS.scala 103:24]
  wire  w_buffer_srst; // @[BFS.scala 103:24]
  wire  w_buffer_valid; // @[BFS.scala 103:24]
  wire  w_buffer_reg_slice_aclk; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_aresetn; // @[BFS.scala 109:34]
  wire [63:0] w_buffer_reg_slice_s_axis_tdata; // @[BFS.scala 109:34]
  wire [7:0] w_buffer_reg_slice_s_axis_tkeep; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tvalid; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tready; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tlast; // @[BFS.scala 109:34]
  wire [63:0] w_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 109:34]
  wire [7:0] w_buffer_reg_slice_m_axis_tkeep; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tready; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tlast; // @[BFS.scala 109:34]
  wire  aw_buffer_reg_slice_aclk; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_aresetn; // @[BFS.scala 112:35]
  wire [63:0] aw_buffer_reg_slice_s_axis_tdata; // @[BFS.scala 112:35]
  wire [7:0] aw_buffer_reg_slice_s_axis_tkeep; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tvalid; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tready; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tlast; // @[BFS.scala 112:35]
  wire [63:0] aw_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 112:35]
  wire [7:0] aw_buffer_reg_slice_m_axis_tkeep; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tready; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tlast; // @[BFS.scala 112:35]
  wire [9:0] block_index = io_xbar_in_bits_tdata[23:14]; // @[BFS.scala 37:8]
  wire [15:0] pipeline_1_out_addr = pipeline_1_m_axis_tdata[27:12]; // @[BFS.scala 69:52]
  wire [11:0] pipeline_1_out_block_index = pipeline_1_m_axis_tdata[11:0]; // @[BFS.scala 70:59]
  wire  _pipeline_1_io_s_axis_tvalid_T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 73:51]
  wire [15:0] pipeline_1_io_s_axis_tdata_hi = {{4'd0}, io_xbar_in_bits_tdata[13:2]}; // @[BFS.scala 41:66 BFS.scala 41:66]
  wire [11:0] pipeline_1_io_s_axis_tdata_lo = {{2'd0}, block_index}; // @[BFS.scala 74:73 BFS.scala 74:73]
  wire [27:0] _pipeline_1_io_s_axis_tdata_T_1 = {pipeline_1_io_s_axis_tdata_hi,pipeline_1_io_s_axis_tdata_lo}; // @[Cat.scala 30:58]
  wire  _buffer_io_wea_T = pipeline_1_m_axis_tvalid; // @[BFS.scala 78:54]
  wire  _buffer_io_wea_T_2 = pipeline_1_m_axis_tvalid & pipeline_1_m_axis_tready; // @[BFS.scala 78:57]
  wire [15:0] _region_counter_doutb_T_1 = region_counter_doutb_forward_m_axis_tvalid ?
    region_counter_doutb_forward_m_axis_tdata : {{7'd0}, region_counter__doutb}; // @[BFS.scala 90:30]
  wire [8:0] region_counter_doutb = _region_counter_doutb_T_1[8:0]; // @[BFS.scala 63:34 BFS.scala 90:24]
  wire [5:0] buffer_io_addra_lo = region_counter_doutb[5:0]; // @[BFS.scala 29:35 BFS.scala 29:35]
  wire [17:0] _buffer_io_addra_T = {pipeline_1_out_block_index,buffer_io_addra_lo}; // @[Cat.scala 30:58]
  wire  _region_counter_dina_0_T = region_counter_doutb == 9'h3f; // @[BFS.scala 33:17]
  wire [8:0] _region_counter_dina_0_T_2 = region_counter_doutb + 9'h1; // @[BFS.scala 33:40]
  wire [8:0] region_counter_dina_0 = region_counter_doutb == 9'h3f ? 9'h0 : _region_counter_dina_0_T_2; // @[BFS.scala 33:8]
  wire  _region_counter_doutb_forward_io_s_axis_tvalid_T_1 = pipeline_1_out_block_index == pipeline_1_io_s_axis_tdata_lo
    ; // @[BFS.scala 88:28]
  wire  _region_counter_doutb_forward_io_s_axis_tvalid_T_2 = _pipeline_1_io_s_axis_tvalid_T &
    _region_counter_doutb_forward_io_s_axis_tvalid_T_1; // @[BFS.scala 87:89]
  reg [1:0] wb_sm; // @[BFS.scala 100:22]
  reg [7:0] count; // @[BFS.scala 101:22]
  reg [9:0] wb_block_index; // @[BFS.scala 104:31]
  wire  _flush_start_T = wb_sm == 2'h0; // @[BFS.scala 105:28]
  wire  flush_start = wb_sm == 2'h0 & io_flush; // @[BFS.scala 105:42]
  reg [7:0] size_b; // @[BFS.scala 106:23]
  reg [63:0] level_base_addr_reg; // @[BFS.scala 107:36]
  wire  wb_start = _buffer_io_wea_T & _region_counter_dina_0_T & _flush_start_T; // @[BFS.scala 108:89]
  wire  _T = wb_sm == 2'h3; // @[BFS.scala 121:20]
  wire [8:0] _GEN_0 = wb_sm == 2'h3 ? region_counter_doutb : {{1'd0}, size_b}; // @[BFS.scala 121:38 BFS.scala 122:12 BFS.scala 106:23]
  wire [8:0] _GEN_1 = wb_start ? 9'h40 : _GEN_0; // @[BFS.scala 119:17 BFS.scala 120:12]
  wire  _T_1 = wb_sm == 2'h2; // @[BFS.scala 129:20]
  wire  _T_2 = wb_block_index != 10'h3ff; // @[BFS.scala 129:55]
  wire [9:0] _wb_block_index_T_1 = wb_block_index + 10'h1; // @[BFS.scala 130:38]
  wire [9:0] _GEN_2 = wb_sm == 2'h2 & wb_block_index != 10'h3ff ? _wb_block_index_T_1 : wb_block_index; // @[BFS.scala 129:72 BFS.scala 130:20 BFS.scala 104:31]
  wire [9:0] _GEN_3 = flush_start ? 10'h0 : _GEN_2; // @[BFS.scala 127:26 BFS.scala 128:20]
  wire [11:0] _GEN_4 = wb_start ? pipeline_1_out_block_index : {{2'd0}, _GEN_3}; // @[BFS.scala 125:17 BFS.scala 126:20]
  wire  _T_6 = wb_sm == 2'h1; // @[BFS.scala 144:20]
  wire  _T_7 = aw_buffer_reg_slice_s_axis_tready; // @[BFS.scala 144:82]
  wire  _T_9 = w_buffer_reg_slice_s_axis_tready; // @[BFS.scala 145:47]
  wire  _T_10 = wb_sm == 2'h1 & aw_buffer_reg_slice_s_axis_tready & _T_9; // @[BFS.scala 144:85]
  wire [1:0] _GEN_6 = io_flush ? 2'h2 : 2'h0; // @[BFS.scala 147:21 BFS.scala 148:15 BFS.scala 150:15]
  wire [1:0] _GEN_7 = count == size_b ? _GEN_6 : 2'h1; // @[BFS.scala 146:27 BFS.scala 153:13]
  wire [1:0] _GEN_8 = _T_2 ? 2'h3 : 2'h0; // @[BFS.scala 156:42 BFS.scala 157:13 BFS.scala 159:13]
  wire [1:0] _GEN_9 = _T_1 ? _GEN_8 : wb_sm; // @[BFS.scala 155:38 BFS.scala 100:22]
  wire [1:0] _GEN_10 = _T_10 ? _GEN_7 : _GEN_9; // @[BFS.scala 145:51]
  wire [7:0] _count_T_1 = count + 8'h1; // @[BFS.scala 167:20]
  wire [15:0] _buffer_io_addrb_T = {block_index,6'h0}; // @[Cat.scala 30:58]
  wire [5:0] buffer_io_addrb_lo_2 = count[5:0]; // @[BFS.scala 29:35 BFS.scala 29:35]
  wire [15:0] _buffer_io_addrb_T_4 = {wb_block_index,buffer_io_addrb_lo_2}; // @[Cat.scala 30:58]
  wire [15:0] _buffer_io_addrb_T_5 = wb_start ? _buffer_io_addrb_T : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_6 = _T ? _buffer_io_addrb_T : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_7 = _T_6 ? _buffer_io_addrb_T_4 : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_8 = _buffer_io_addrb_T_5 | _buffer_io_addrb_T_6; // @[Mux.scala 27:72]
  wire [11:0] _region_counter_io_addra_T_1 = _T_6 ? {{2'd0}, wb_block_index} : pipeline_1_out_block_index; // @[BFS.scala 180:33]
  wire [11:0] _region_counter_io_addrb_T_4 = _T_6 ? pipeline_1_out_block_index : {{2'd0}, block_index}; // @[Mux.scala 98:16]
  wire [11:0] _region_counter_io_addrb_T_5 = flush_start ? 12'h0 : _region_counter_io_addrb_T_4; // @[Mux.scala 98:16]
  wire [11:0] _region_counter_io_addrb_T_6 = _T_1 ? {{2'd0}, _wb_block_index_T_1} : _region_counter_io_addrb_T_5; // @[Mux.scala 98:16]
  wire [11:0] aw_buffer_reg_slice_io_s_axis_tdata_lo = buffer_io_doutb[43:32]; // @[BFS.scala 45:43]
  wire [23:0] _aw_buffer_reg_slice_io_s_axis_tdata_T_1 = {wb_block_index,2'h0,aw_buffer_reg_slice_io_s_axis_tdata_lo}; // @[Cat.scala 30:58]
  wire [25:0] _aw_buffer_reg_slice_io_s_axis_tdata_T_2 = {_aw_buffer_reg_slice_io_s_axis_tdata_T_1, 2'h0}; // @[BFS.scala 45:53]
  wire [59:0] alignment_addr = aw_buffer_dout[63:4]; // @[BFS.scala 196:41]
  wire [4:0] io_axi_ddr_aw_bits_awid_lo = aw_buffer_data_count[4:0]; // @[BFS.scala 199:76 BFS.scala 199:76]
  wire [3:0] alignment_offset = {w_buffer_dout[33:32], 2'h0}; // @[BFS.scala 213:52]
  wire [7:0] _io_axi_ddr_w_bits_wdata_T_1 = 4'h8 * alignment_offset; // @[BFS.scala 214:84]
  wire [127:0] _io_axi_ddr_w_bits_wdata_WIRE = {{96'd0}, w_buffer_dout[31:0]}; // @[BFS.scala 214:62 BFS.scala 214:62]
  wire [382:0] _GEN_17 = {{255'd0}, _io_axi_ddr_w_bits_wdata_WIRE}; // @[BFS.scala 214:76]
  wire [382:0] _io_axi_ddr_w_bits_wdata_T_2 = _GEN_17 << _io_axi_ddr_w_bits_wdata_T_1; // @[BFS.scala 214:76]
  wire [30:0] _io_axi_ddr_w_bits_wstrb_T = 31'hf << alignment_offset; // @[BFS.scala 217:42]
  URAM_cluster buffer ( // @[BFS.scala 25:22]
    .io_addra(buffer_io_addra),
    .io_clka(buffer_io_clka),
    .io_dina(buffer_io_dina),
    .io_wea(buffer_io_wea),
    .io_addrb(buffer_io_addrb),
    .io_clkb(buffer_io_clkb),
    .io_doutb(buffer_io_doutb)
  );
  region_counter region_counter_ ( // @[BFS.scala 26:30]
    .addra(region_counter__addra),
    .clka(region_counter__clka),
    .dina(region_counter__dina),
    .ena(region_counter__ena),
    .wea(region_counter__wea),
    .addrb(region_counter__addrb),
    .clkb(region_counter__clkb),
    .doutb(region_counter__doutb),
    .enb(region_counter__enb)
  );
  region_counter_doutb_forward_reg_slice region_counter_doutb_forward ( // @[BFS.scala 60:44]
    .aclk(region_counter_doutb_forward_aclk),
    .aresetn(region_counter_doutb_forward_aresetn),
    .s_axis_tdata(region_counter_doutb_forward_s_axis_tdata),
    .s_axis_tkeep(region_counter_doutb_forward_s_axis_tkeep),
    .s_axis_tvalid(region_counter_doutb_forward_s_axis_tvalid),
    .s_axis_tready(region_counter_doutb_forward_s_axis_tready),
    .s_axis_tlast(region_counter_doutb_forward_s_axis_tlast),
    .m_axis_tdata(region_counter_doutb_forward_m_axis_tdata),
    .m_axis_tkeep(region_counter_doutb_forward_m_axis_tkeep),
    .m_axis_tvalid(region_counter_doutb_forward_m_axis_tvalid),
    .m_axis_tready(region_counter_doutb_forward_m_axis_tready),
    .m_axis_tlast(region_counter_doutb_forward_m_axis_tlast)
  );
  WB_engine_in_reg_slice pipeline_1 ( // @[BFS.scala 64:26]
    .aclk(pipeline_1_aclk),
    .aresetn(pipeline_1_aresetn),
    .s_axis_tdata(pipeline_1_s_axis_tdata),
    .s_axis_tkeep(pipeline_1_s_axis_tkeep),
    .s_axis_tvalid(pipeline_1_s_axis_tvalid),
    .s_axis_tready(pipeline_1_s_axis_tready),
    .s_axis_tlast(pipeline_1_s_axis_tlast),
    .m_axis_tdata(pipeline_1_m_axis_tdata),
    .m_axis_tkeep(pipeline_1_m_axis_tkeep),
    .m_axis_tvalid(pipeline_1_m_axis_tvalid),
    .m_axis_tready(pipeline_1_m_axis_tready),
    .m_axis_tlast(pipeline_1_m_axis_tlast)
  );
  addr_fifo aw_buffer ( // @[BFS.scala 102:25]
    .full(aw_buffer_full),
    .din(aw_buffer_din),
    .wr_en(aw_buffer_wr_en),
    .empty(aw_buffer_empty),
    .dout(aw_buffer_dout),
    .rd_en(aw_buffer_rd_en),
    .data_count(aw_buffer_data_count),
    .clk(aw_buffer_clk),
    .srst(aw_buffer_srst),
    .valid(aw_buffer_valid)
  );
  level_fifo w_buffer ( // @[BFS.scala 103:24]
    .full(w_buffer_full),
    .din(w_buffer_din),
    .wr_en(w_buffer_wr_en),
    .empty(w_buffer_empty),
    .dout(w_buffer_dout),
    .rd_en(w_buffer_rd_en),
    .data_count(w_buffer_data_count),
    .clk(w_buffer_clk),
    .srst(w_buffer_srst),
    .valid(w_buffer_valid)
  );
  w_buffer_reg_slice w_buffer_reg_slice ( // @[BFS.scala 109:34]
    .aclk(w_buffer_reg_slice_aclk),
    .aresetn(w_buffer_reg_slice_aresetn),
    .s_axis_tdata(w_buffer_reg_slice_s_axis_tdata),
    .s_axis_tkeep(w_buffer_reg_slice_s_axis_tkeep),
    .s_axis_tvalid(w_buffer_reg_slice_s_axis_tvalid),
    .s_axis_tready(w_buffer_reg_slice_s_axis_tready),
    .s_axis_tlast(w_buffer_reg_slice_s_axis_tlast),
    .m_axis_tdata(w_buffer_reg_slice_m_axis_tdata),
    .m_axis_tkeep(w_buffer_reg_slice_m_axis_tkeep),
    .m_axis_tvalid(w_buffer_reg_slice_m_axis_tvalid),
    .m_axis_tready(w_buffer_reg_slice_m_axis_tready),
    .m_axis_tlast(w_buffer_reg_slice_m_axis_tlast)
  );
  aw_buffer_reg_slice aw_buffer_reg_slice ( // @[BFS.scala 112:35]
    .aclk(aw_buffer_reg_slice_aclk),
    .aresetn(aw_buffer_reg_slice_aresetn),
    .s_axis_tdata(aw_buffer_reg_slice_s_axis_tdata),
    .s_axis_tkeep(aw_buffer_reg_slice_s_axis_tkeep),
    .s_axis_tvalid(aw_buffer_reg_slice_s_axis_tvalid),
    .s_axis_tready(aw_buffer_reg_slice_s_axis_tready),
    .s_axis_tlast(aw_buffer_reg_slice_s_axis_tlast),
    .m_axis_tdata(aw_buffer_reg_slice_m_axis_tdata),
    .m_axis_tkeep(aw_buffer_reg_slice_m_axis_tkeep),
    .m_axis_tvalid(aw_buffer_reg_slice_m_axis_tvalid),
    .m_axis_tready(aw_buffer_reg_slice_m_axis_tready),
    .m_axis_tlast(aw_buffer_reg_slice_m_axis_tlast)
  );
  assign io_axi_ddr_aw_valid = aw_buffer_valid; // @[BFS.scala 203:23]
  assign io_axi_ddr_aw_bits_awaddr = {alignment_addr,4'h0}; // @[Cat.scala 30:58]
  assign io_axi_ddr_aw_bits_awid = {1'h1,io_axi_ddr_aw_bits_awid_lo}; // @[Cat.scala 30:58]
  assign io_axi_ddr_w_valid = w_buffer_valid; // @[BFS.scala 216:22]
  assign io_axi_ddr_w_bits_wdata = _io_axi_ddr_w_bits_wdata_T_2[127:0]; // @[BFS.scala 214:27]
  assign io_axi_ddr_w_bits_wstrb = _io_axi_ddr_w_bits_wstrb_T[15:0]; // @[BFS.scala 217:27]
  assign io_xbar_in_ready = pipeline_1_s_axis_tready; // @[BFS.scala 75:20]
  assign io_end = _T_1 & wb_block_index == 10'h3ff; // @[BFS.scala 221:36]
  assign buffer_io_addra = _buffer_io_addra_T[15:0]; // @[BFS.scala 79:19]
  assign buffer_io_clka = clock; // @[BFS.scala 81:33]
  assign buffer_io_dina = {pipeline_1_out_addr,io_level}; // @[Cat.scala 30:58]
  assign buffer_io_wea = pipeline_1_m_axis_tvalid & pipeline_1_m_axis_tready; // @[BFS.scala 78:57]
  assign buffer_io_addrb = _buffer_io_addrb_T_8 | _buffer_io_addrb_T_7; // @[Mux.scala 27:72]
  assign buffer_io_clkb = clock; // @[BFS.scala 178:33]
  assign region_counter__addra = _region_counter_io_addra_T_1[9:0]; // @[BFS.scala 180:27]
  assign region_counter__clka = clock; // @[BFS.scala 54:41]
  assign region_counter__dina = _T_6 ? 9'h0 : region_counter_dina_0; // @[BFS.scala 182:32]
  assign region_counter__ena = 1'h1; // @[BFS.scala 55:25]
  assign region_counter__wea = _T_6 | _buffer_io_wea_T_2; // @[BFS.scala 181:31]
  assign region_counter__addrb = _region_counter_io_addrb_T_6[9:0]; // @[BFS.scala 183:27]
  assign region_counter__clkb = clock; // @[BFS.scala 53:41]
  assign region_counter__enb = 1'h1; // @[BFS.scala 56:25]
  assign region_counter_doutb_forward_aclk = clock; // @[BFS.scala 61:55]
  assign region_counter_doutb_forward_aresetn = ~reset; // @[BFS.scala 62:46]
  assign region_counter_doutb_forward_s_axis_tdata = {{7'd0}, region_counter_dina_0}; // @[BFS.scala 33:8]
  assign region_counter_doutb_forward_s_axis_tkeep = 2'h0;
  assign region_counter_doutb_forward_s_axis_tvalid = _region_counter_doutb_forward_io_s_axis_tvalid_T_2 &
    _buffer_io_wea_T_2; // @[BFS.scala 88:55]
  assign region_counter_doutb_forward_s_axis_tlast = 1'h0;
  assign region_counter_doutb_forward_m_axis_tready = wb_sm == 2'h0; // @[BFS.scala 116:58]
  assign pipeline_1_aclk = clock; // @[BFS.scala 71:37]
  assign pipeline_1_aresetn = ~reset; // @[BFS.scala 72:28]
  assign pipeline_1_s_axis_tdata = {{4'd0}, _pipeline_1_io_s_axis_tdata_T_1}; // @[Cat.scala 30:58]
  assign pipeline_1_s_axis_tkeep = 4'h0;
  assign pipeline_1_s_axis_tvalid = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 73:51]
  assign pipeline_1_s_axis_tlast = 1'h0;
  assign pipeline_1_m_axis_tready = wb_sm == 2'h0; // @[BFS.scala 115:40]
  assign aw_buffer_din = aw_buffer_reg_slice_m_axis_tdata + level_base_addr_reg; // @[BFS.scala 195:59]
  assign aw_buffer_wr_en = aw_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 194:22]
  assign aw_buffer_rd_en = io_axi_ddr_aw_ready; // @[BFS.scala 204:22]
  assign aw_buffer_clk = clock; // @[BFS.scala 192:35]
  assign aw_buffer_srst = reset; // @[BFS.scala 193:36]
  assign w_buffer_din = w_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 212:19]
  assign w_buffer_wr_en = w_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 211:21]
  assign w_buffer_rd_en = io_axi_ddr_w_ready; // @[BFS.scala 218:21]
  assign w_buffer_clk = clock; // @[BFS.scala 209:34]
  assign w_buffer_srst = reset; // @[BFS.scala 210:35]
  assign w_buffer_reg_slice_aclk = clock; // @[BFS.scala 110:45]
  assign w_buffer_reg_slice_aresetn = ~reset; // @[BFS.scala 111:36]
  assign w_buffer_reg_slice_s_axis_tdata = {{30'd0}, buffer_io_doutb[33:0]}; // @[BFS.scala 206:56]
  assign w_buffer_reg_slice_s_axis_tkeep = 8'h0;
  assign w_buffer_reg_slice_s_axis_tvalid = _T_6 & _T_7; // @[BFS.scala 207:64]
  assign w_buffer_reg_slice_s_axis_tlast = 1'h0;
  assign w_buffer_reg_slice_m_axis_tready = ~w_buffer_full; // @[util.scala 219:13]
  assign aw_buffer_reg_slice_aclk = clock; // @[BFS.scala 113:46]
  assign aw_buffer_reg_slice_aresetn = ~reset; // @[BFS.scala 114:37]
  assign aw_buffer_reg_slice_s_axis_tdata = {{38'd0}, _aw_buffer_reg_slice_io_s_axis_tdata_T_2}; // @[BFS.scala 45:53]
  assign aw_buffer_reg_slice_s_axis_tkeep = 8'h0;
  assign aw_buffer_reg_slice_s_axis_tvalid = _T_6 & _T_9; // @[BFS.scala 190:65]
  assign aw_buffer_reg_slice_s_axis_tlast = 1'h0;
  assign aw_buffer_reg_slice_m_axis_tready = ~aw_buffer_full; // @[util.scala 219:13]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 100:22]
      wb_sm <= 2'h0; // @[BFS.scala 100:22]
    end else if (flush_start) begin // @[BFS.scala 134:20]
      wb_sm <= 2'h3; // @[BFS.scala 135:11]
    end else if (_T) begin // @[BFS.scala 136:38]
      if (region_counter_doutb == 9'h0) begin // @[BFS.scala 137:39]
        wb_sm <= 2'h2; // @[BFS.scala 138:13]
      end else begin
        wb_sm <= 2'h1; // @[BFS.scala 140:13]
      end
    end else if (wb_start) begin // @[BFS.scala 142:23]
      wb_sm <= 2'h1; // @[BFS.scala 143:11]
    end else begin
      wb_sm <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 101:22]
      count <= 8'h0; // @[BFS.scala 101:22]
    end else if (_flush_start_T | _T_1) begin // @[BFS.scala 163:53]
      count <= 8'h1; // @[BFS.scala 164:11]
    end else if (_T_10) begin // @[BFS.scala 166:50]
      count <= _count_T_1; // @[BFS.scala 167:11]
    end
    if (reset) begin // @[BFS.scala 104:31]
      wb_block_index <= 10'h0; // @[BFS.scala 104:31]
    end else begin
      wb_block_index <= _GEN_4[9:0];
    end
    if (reset) begin // @[BFS.scala 106:23]
      size_b <= 8'h0; // @[BFS.scala 106:23]
    end else begin
      size_b <= _GEN_1[7:0];
    end
    if (reset) begin // @[BFS.scala 107:36]
      level_base_addr_reg <= 64'h0; // @[BFS.scala 107:36]
    end else begin
      level_base_addr_reg <= io_level_base_addr; // @[BFS.scala 117:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_sm = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  wb_block_index = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  size_b = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  level_base_addr_reg = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WB_engine_1(
  input          clock,
  input          reset,
  input          io_axi_ddr_aw_ready,
  output         io_axi_ddr_aw_valid,
  output [63:0]  io_axi_ddr_aw_bits_awaddr,
  output [5:0]   io_axi_ddr_aw_bits_awid,
  input          io_axi_ddr_w_ready,
  output         io_axi_ddr_w_valid,
  output [127:0] io_axi_ddr_w_bits_wdata,
  output [15:0]  io_axi_ddr_w_bits_wstrb,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [31:0]  io_xbar_in_bits_tdata,
  input  [63:0]  io_level_base_addr,
  input  [31:0]  io_level,
  output         io_end,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] buffer_io_addra; // @[BFS.scala 25:22]
  wire  buffer_io_clka; // @[BFS.scala 25:22]
  wire [47:0] buffer_io_dina; // @[BFS.scala 25:22]
  wire  buffer_io_wea; // @[BFS.scala 25:22]
  wire [15:0] buffer_io_addrb; // @[BFS.scala 25:22]
  wire  buffer_io_clkb; // @[BFS.scala 25:22]
  wire [47:0] buffer_io_doutb; // @[BFS.scala 25:22]
  wire [9:0] region_counter__addra; // @[BFS.scala 26:30]
  wire  region_counter__clka; // @[BFS.scala 26:30]
  wire [8:0] region_counter__dina; // @[BFS.scala 26:30]
  wire  region_counter__ena; // @[BFS.scala 26:30]
  wire  region_counter__wea; // @[BFS.scala 26:30]
  wire [9:0] region_counter__addrb; // @[BFS.scala 26:30]
  wire  region_counter__clkb; // @[BFS.scala 26:30]
  wire [8:0] region_counter__doutb; // @[BFS.scala 26:30]
  wire  region_counter__enb; // @[BFS.scala 26:30]
  wire  region_counter_doutb_forward_aclk; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_aresetn; // @[BFS.scala 60:44]
  wire [15:0] region_counter_doutb_forward_s_axis_tdata; // @[BFS.scala 60:44]
  wire [1:0] region_counter_doutb_forward_s_axis_tkeep; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tvalid; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tready; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tlast; // @[BFS.scala 60:44]
  wire [15:0] region_counter_doutb_forward_m_axis_tdata; // @[BFS.scala 60:44]
  wire [1:0] region_counter_doutb_forward_m_axis_tkeep; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tvalid; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tready; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tlast; // @[BFS.scala 60:44]
  wire  pipeline_1_aclk; // @[BFS.scala 64:26]
  wire  pipeline_1_aresetn; // @[BFS.scala 64:26]
  wire [31:0] pipeline_1_s_axis_tdata; // @[BFS.scala 64:26]
  wire [3:0] pipeline_1_s_axis_tkeep; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tvalid; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tready; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tlast; // @[BFS.scala 64:26]
  wire [31:0] pipeline_1_m_axis_tdata; // @[BFS.scala 64:26]
  wire [3:0] pipeline_1_m_axis_tkeep; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tvalid; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tready; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tlast; // @[BFS.scala 64:26]
  wire  aw_buffer_full; // @[BFS.scala 102:25]
  wire [63:0] aw_buffer_din; // @[BFS.scala 102:25]
  wire  aw_buffer_wr_en; // @[BFS.scala 102:25]
  wire  aw_buffer_empty; // @[BFS.scala 102:25]
  wire [63:0] aw_buffer_dout; // @[BFS.scala 102:25]
  wire  aw_buffer_rd_en; // @[BFS.scala 102:25]
  wire [5:0] aw_buffer_data_count; // @[BFS.scala 102:25]
  wire  aw_buffer_clk; // @[BFS.scala 102:25]
  wire  aw_buffer_srst; // @[BFS.scala 102:25]
  wire  aw_buffer_valid; // @[BFS.scala 102:25]
  wire  w_buffer_full; // @[BFS.scala 103:24]
  wire [63:0] w_buffer_din; // @[BFS.scala 103:24]
  wire  w_buffer_wr_en; // @[BFS.scala 103:24]
  wire  w_buffer_empty; // @[BFS.scala 103:24]
  wire [63:0] w_buffer_dout; // @[BFS.scala 103:24]
  wire  w_buffer_rd_en; // @[BFS.scala 103:24]
  wire [5:0] w_buffer_data_count; // @[BFS.scala 103:24]
  wire  w_buffer_clk; // @[BFS.scala 103:24]
  wire  w_buffer_srst; // @[BFS.scala 103:24]
  wire  w_buffer_valid; // @[BFS.scala 103:24]
  wire  w_buffer_reg_slice_aclk; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_aresetn; // @[BFS.scala 109:34]
  wire [63:0] w_buffer_reg_slice_s_axis_tdata; // @[BFS.scala 109:34]
  wire [7:0] w_buffer_reg_slice_s_axis_tkeep; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tvalid; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tready; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tlast; // @[BFS.scala 109:34]
  wire [63:0] w_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 109:34]
  wire [7:0] w_buffer_reg_slice_m_axis_tkeep; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tready; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tlast; // @[BFS.scala 109:34]
  wire  aw_buffer_reg_slice_aclk; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_aresetn; // @[BFS.scala 112:35]
  wire [63:0] aw_buffer_reg_slice_s_axis_tdata; // @[BFS.scala 112:35]
  wire [7:0] aw_buffer_reg_slice_s_axis_tkeep; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tvalid; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tready; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tlast; // @[BFS.scala 112:35]
  wire [63:0] aw_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 112:35]
  wire [7:0] aw_buffer_reg_slice_m_axis_tkeep; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tready; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tlast; // @[BFS.scala 112:35]
  wire [9:0] block_index = io_xbar_in_bits_tdata[23:14]; // @[BFS.scala 37:8]
  wire [15:0] pipeline_1_out_addr = pipeline_1_m_axis_tdata[27:12]; // @[BFS.scala 69:52]
  wire [11:0] pipeline_1_out_block_index = pipeline_1_m_axis_tdata[11:0]; // @[BFS.scala 70:59]
  wire  _pipeline_1_io_s_axis_tvalid_T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 73:51]
  wire [15:0] pipeline_1_io_s_axis_tdata_hi = {{4'd0}, io_xbar_in_bits_tdata[13:2]}; // @[BFS.scala 41:66 BFS.scala 41:66]
  wire [11:0] pipeline_1_io_s_axis_tdata_lo = {{2'd0}, block_index}; // @[BFS.scala 74:73 BFS.scala 74:73]
  wire [27:0] _pipeline_1_io_s_axis_tdata_T_1 = {pipeline_1_io_s_axis_tdata_hi,pipeline_1_io_s_axis_tdata_lo}; // @[Cat.scala 30:58]
  wire  _buffer_io_wea_T = pipeline_1_m_axis_tvalid; // @[BFS.scala 78:54]
  wire  _buffer_io_wea_T_2 = pipeline_1_m_axis_tvalid & pipeline_1_m_axis_tready; // @[BFS.scala 78:57]
  wire [15:0] _region_counter_doutb_T_1 = region_counter_doutb_forward_m_axis_tvalid ?
    region_counter_doutb_forward_m_axis_tdata : {{7'd0}, region_counter__doutb}; // @[BFS.scala 90:30]
  wire [8:0] region_counter_doutb = _region_counter_doutb_T_1[8:0]; // @[BFS.scala 63:34 BFS.scala 90:24]
  wire [5:0] buffer_io_addra_lo = region_counter_doutb[5:0]; // @[BFS.scala 29:35 BFS.scala 29:35]
  wire [17:0] _buffer_io_addra_T = {pipeline_1_out_block_index,buffer_io_addra_lo}; // @[Cat.scala 30:58]
  wire  _region_counter_dina_0_T = region_counter_doutb == 9'h3f; // @[BFS.scala 33:17]
  wire [8:0] _region_counter_dina_0_T_2 = region_counter_doutb + 9'h1; // @[BFS.scala 33:40]
  wire [8:0] region_counter_dina_0 = region_counter_doutb == 9'h3f ? 9'h0 : _region_counter_dina_0_T_2; // @[BFS.scala 33:8]
  wire  _region_counter_doutb_forward_io_s_axis_tvalid_T_1 = pipeline_1_out_block_index == pipeline_1_io_s_axis_tdata_lo
    ; // @[BFS.scala 88:28]
  wire  _region_counter_doutb_forward_io_s_axis_tvalid_T_2 = _pipeline_1_io_s_axis_tvalid_T &
    _region_counter_doutb_forward_io_s_axis_tvalid_T_1; // @[BFS.scala 87:89]
  reg [1:0] wb_sm; // @[BFS.scala 100:22]
  reg [7:0] count; // @[BFS.scala 101:22]
  reg [9:0] wb_block_index; // @[BFS.scala 104:31]
  wire  _flush_start_T = wb_sm == 2'h0; // @[BFS.scala 105:28]
  wire  flush_start = wb_sm == 2'h0 & io_flush; // @[BFS.scala 105:42]
  reg [7:0] size_b; // @[BFS.scala 106:23]
  reg [63:0] level_base_addr_reg; // @[BFS.scala 107:36]
  wire  wb_start = _buffer_io_wea_T & _region_counter_dina_0_T & _flush_start_T; // @[BFS.scala 108:89]
  wire  _T = wb_sm == 2'h3; // @[BFS.scala 121:20]
  wire [8:0] _GEN_0 = wb_sm == 2'h3 ? region_counter_doutb : {{1'd0}, size_b}; // @[BFS.scala 121:38 BFS.scala 122:12 BFS.scala 106:23]
  wire [8:0] _GEN_1 = wb_start ? 9'h40 : _GEN_0; // @[BFS.scala 119:17 BFS.scala 120:12]
  wire  _T_1 = wb_sm == 2'h2; // @[BFS.scala 129:20]
  wire  _T_2 = wb_block_index != 10'h3ff; // @[BFS.scala 129:55]
  wire [9:0] _wb_block_index_T_1 = wb_block_index + 10'h1; // @[BFS.scala 130:38]
  wire [9:0] _GEN_2 = wb_sm == 2'h2 & wb_block_index != 10'h3ff ? _wb_block_index_T_1 : wb_block_index; // @[BFS.scala 129:72 BFS.scala 130:20 BFS.scala 104:31]
  wire [9:0] _GEN_3 = flush_start ? 10'h0 : _GEN_2; // @[BFS.scala 127:26 BFS.scala 128:20]
  wire [11:0] _GEN_4 = wb_start ? pipeline_1_out_block_index : {{2'd0}, _GEN_3}; // @[BFS.scala 125:17 BFS.scala 126:20]
  wire  _T_6 = wb_sm == 2'h1; // @[BFS.scala 144:20]
  wire  _T_7 = aw_buffer_reg_slice_s_axis_tready; // @[BFS.scala 144:82]
  wire  _T_9 = w_buffer_reg_slice_s_axis_tready; // @[BFS.scala 145:47]
  wire  _T_10 = wb_sm == 2'h1 & aw_buffer_reg_slice_s_axis_tready & _T_9; // @[BFS.scala 144:85]
  wire [1:0] _GEN_6 = io_flush ? 2'h2 : 2'h0; // @[BFS.scala 147:21 BFS.scala 148:15 BFS.scala 150:15]
  wire [1:0] _GEN_7 = count == size_b ? _GEN_6 : 2'h1; // @[BFS.scala 146:27 BFS.scala 153:13]
  wire [1:0] _GEN_8 = _T_2 ? 2'h3 : 2'h0; // @[BFS.scala 156:42 BFS.scala 157:13 BFS.scala 159:13]
  wire [1:0] _GEN_9 = _T_1 ? _GEN_8 : wb_sm; // @[BFS.scala 155:38 BFS.scala 100:22]
  wire [1:0] _GEN_10 = _T_10 ? _GEN_7 : _GEN_9; // @[BFS.scala 145:51]
  wire [7:0] _count_T_1 = count + 8'h1; // @[BFS.scala 167:20]
  wire [15:0] _buffer_io_addrb_T = {block_index,6'h0}; // @[Cat.scala 30:58]
  wire [5:0] buffer_io_addrb_lo_2 = count[5:0]; // @[BFS.scala 29:35 BFS.scala 29:35]
  wire [15:0] _buffer_io_addrb_T_4 = {wb_block_index,buffer_io_addrb_lo_2}; // @[Cat.scala 30:58]
  wire [15:0] _buffer_io_addrb_T_5 = wb_start ? _buffer_io_addrb_T : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_6 = _T ? _buffer_io_addrb_T : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_7 = _T_6 ? _buffer_io_addrb_T_4 : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_8 = _buffer_io_addrb_T_5 | _buffer_io_addrb_T_6; // @[Mux.scala 27:72]
  wire [11:0] _region_counter_io_addra_T_1 = _T_6 ? {{2'd0}, wb_block_index} : pipeline_1_out_block_index; // @[BFS.scala 180:33]
  wire [11:0] _region_counter_io_addrb_T_4 = _T_6 ? pipeline_1_out_block_index : {{2'd0}, block_index}; // @[Mux.scala 98:16]
  wire [11:0] _region_counter_io_addrb_T_5 = flush_start ? 12'h0 : _region_counter_io_addrb_T_4; // @[Mux.scala 98:16]
  wire [11:0] _region_counter_io_addrb_T_6 = _T_1 ? {{2'd0}, _wb_block_index_T_1} : _region_counter_io_addrb_T_5; // @[Mux.scala 98:16]
  wire [11:0] aw_buffer_reg_slice_io_s_axis_tdata_lo = buffer_io_doutb[43:32]; // @[BFS.scala 45:43]
  wire [23:0] _aw_buffer_reg_slice_io_s_axis_tdata_T_1 = {wb_block_index,2'h1,aw_buffer_reg_slice_io_s_axis_tdata_lo}; // @[Cat.scala 30:58]
  wire [25:0] _aw_buffer_reg_slice_io_s_axis_tdata_T_2 = {_aw_buffer_reg_slice_io_s_axis_tdata_T_1, 2'h0}; // @[BFS.scala 45:53]
  wire [59:0] alignment_addr = aw_buffer_dout[63:4]; // @[BFS.scala 196:41]
  wire [4:0] io_axi_ddr_aw_bits_awid_lo = aw_buffer_data_count[4:0]; // @[BFS.scala 199:76 BFS.scala 199:76]
  wire [3:0] alignment_offset = {w_buffer_dout[33:32], 2'h0}; // @[BFS.scala 213:52]
  wire [7:0] _io_axi_ddr_w_bits_wdata_T_1 = 4'h8 * alignment_offset; // @[BFS.scala 214:84]
  wire [127:0] _io_axi_ddr_w_bits_wdata_WIRE = {{96'd0}, w_buffer_dout[31:0]}; // @[BFS.scala 214:62 BFS.scala 214:62]
  wire [382:0] _GEN_17 = {{255'd0}, _io_axi_ddr_w_bits_wdata_WIRE}; // @[BFS.scala 214:76]
  wire [382:0] _io_axi_ddr_w_bits_wdata_T_2 = _GEN_17 << _io_axi_ddr_w_bits_wdata_T_1; // @[BFS.scala 214:76]
  wire [30:0] _io_axi_ddr_w_bits_wstrb_T = 31'hf << alignment_offset; // @[BFS.scala 217:42]
  URAM_cluster buffer ( // @[BFS.scala 25:22]
    .io_addra(buffer_io_addra),
    .io_clka(buffer_io_clka),
    .io_dina(buffer_io_dina),
    .io_wea(buffer_io_wea),
    .io_addrb(buffer_io_addrb),
    .io_clkb(buffer_io_clkb),
    .io_doutb(buffer_io_doutb)
  );
  region_counter region_counter_ ( // @[BFS.scala 26:30]
    .addra(region_counter__addra),
    .clka(region_counter__clka),
    .dina(region_counter__dina),
    .ena(region_counter__ena),
    .wea(region_counter__wea),
    .addrb(region_counter__addrb),
    .clkb(region_counter__clkb),
    .doutb(region_counter__doutb),
    .enb(region_counter__enb)
  );
  region_counter_doutb_forward_reg_slice region_counter_doutb_forward ( // @[BFS.scala 60:44]
    .aclk(region_counter_doutb_forward_aclk),
    .aresetn(region_counter_doutb_forward_aresetn),
    .s_axis_tdata(region_counter_doutb_forward_s_axis_tdata),
    .s_axis_tkeep(region_counter_doutb_forward_s_axis_tkeep),
    .s_axis_tvalid(region_counter_doutb_forward_s_axis_tvalid),
    .s_axis_tready(region_counter_doutb_forward_s_axis_tready),
    .s_axis_tlast(region_counter_doutb_forward_s_axis_tlast),
    .m_axis_tdata(region_counter_doutb_forward_m_axis_tdata),
    .m_axis_tkeep(region_counter_doutb_forward_m_axis_tkeep),
    .m_axis_tvalid(region_counter_doutb_forward_m_axis_tvalid),
    .m_axis_tready(region_counter_doutb_forward_m_axis_tready),
    .m_axis_tlast(region_counter_doutb_forward_m_axis_tlast)
  );
  WB_engine_in_reg_slice pipeline_1 ( // @[BFS.scala 64:26]
    .aclk(pipeline_1_aclk),
    .aresetn(pipeline_1_aresetn),
    .s_axis_tdata(pipeline_1_s_axis_tdata),
    .s_axis_tkeep(pipeline_1_s_axis_tkeep),
    .s_axis_tvalid(pipeline_1_s_axis_tvalid),
    .s_axis_tready(pipeline_1_s_axis_tready),
    .s_axis_tlast(pipeline_1_s_axis_tlast),
    .m_axis_tdata(pipeline_1_m_axis_tdata),
    .m_axis_tkeep(pipeline_1_m_axis_tkeep),
    .m_axis_tvalid(pipeline_1_m_axis_tvalid),
    .m_axis_tready(pipeline_1_m_axis_tready),
    .m_axis_tlast(pipeline_1_m_axis_tlast)
  );
  addr_fifo aw_buffer ( // @[BFS.scala 102:25]
    .full(aw_buffer_full),
    .din(aw_buffer_din),
    .wr_en(aw_buffer_wr_en),
    .empty(aw_buffer_empty),
    .dout(aw_buffer_dout),
    .rd_en(aw_buffer_rd_en),
    .data_count(aw_buffer_data_count),
    .clk(aw_buffer_clk),
    .srst(aw_buffer_srst),
    .valid(aw_buffer_valid)
  );
  level_fifo w_buffer ( // @[BFS.scala 103:24]
    .full(w_buffer_full),
    .din(w_buffer_din),
    .wr_en(w_buffer_wr_en),
    .empty(w_buffer_empty),
    .dout(w_buffer_dout),
    .rd_en(w_buffer_rd_en),
    .data_count(w_buffer_data_count),
    .clk(w_buffer_clk),
    .srst(w_buffer_srst),
    .valid(w_buffer_valid)
  );
  w_buffer_reg_slice w_buffer_reg_slice ( // @[BFS.scala 109:34]
    .aclk(w_buffer_reg_slice_aclk),
    .aresetn(w_buffer_reg_slice_aresetn),
    .s_axis_tdata(w_buffer_reg_slice_s_axis_tdata),
    .s_axis_tkeep(w_buffer_reg_slice_s_axis_tkeep),
    .s_axis_tvalid(w_buffer_reg_slice_s_axis_tvalid),
    .s_axis_tready(w_buffer_reg_slice_s_axis_tready),
    .s_axis_tlast(w_buffer_reg_slice_s_axis_tlast),
    .m_axis_tdata(w_buffer_reg_slice_m_axis_tdata),
    .m_axis_tkeep(w_buffer_reg_slice_m_axis_tkeep),
    .m_axis_tvalid(w_buffer_reg_slice_m_axis_tvalid),
    .m_axis_tready(w_buffer_reg_slice_m_axis_tready),
    .m_axis_tlast(w_buffer_reg_slice_m_axis_tlast)
  );
  aw_buffer_reg_slice aw_buffer_reg_slice ( // @[BFS.scala 112:35]
    .aclk(aw_buffer_reg_slice_aclk),
    .aresetn(aw_buffer_reg_slice_aresetn),
    .s_axis_tdata(aw_buffer_reg_slice_s_axis_tdata),
    .s_axis_tkeep(aw_buffer_reg_slice_s_axis_tkeep),
    .s_axis_tvalid(aw_buffer_reg_slice_s_axis_tvalid),
    .s_axis_tready(aw_buffer_reg_slice_s_axis_tready),
    .s_axis_tlast(aw_buffer_reg_slice_s_axis_tlast),
    .m_axis_tdata(aw_buffer_reg_slice_m_axis_tdata),
    .m_axis_tkeep(aw_buffer_reg_slice_m_axis_tkeep),
    .m_axis_tvalid(aw_buffer_reg_slice_m_axis_tvalid),
    .m_axis_tready(aw_buffer_reg_slice_m_axis_tready),
    .m_axis_tlast(aw_buffer_reg_slice_m_axis_tlast)
  );
  assign io_axi_ddr_aw_valid = aw_buffer_valid; // @[BFS.scala 203:23]
  assign io_axi_ddr_aw_bits_awaddr = {alignment_addr,4'h0}; // @[Cat.scala 30:58]
  assign io_axi_ddr_aw_bits_awid = {1'h1,io_axi_ddr_aw_bits_awid_lo}; // @[Cat.scala 30:58]
  assign io_axi_ddr_w_valid = w_buffer_valid; // @[BFS.scala 216:22]
  assign io_axi_ddr_w_bits_wdata = _io_axi_ddr_w_bits_wdata_T_2[127:0]; // @[BFS.scala 214:27]
  assign io_axi_ddr_w_bits_wstrb = _io_axi_ddr_w_bits_wstrb_T[15:0]; // @[BFS.scala 217:27]
  assign io_xbar_in_ready = pipeline_1_s_axis_tready; // @[BFS.scala 75:20]
  assign io_end = _T_1 & wb_block_index == 10'h3ff; // @[BFS.scala 221:36]
  assign buffer_io_addra = _buffer_io_addra_T[15:0]; // @[BFS.scala 79:19]
  assign buffer_io_clka = clock; // @[BFS.scala 81:33]
  assign buffer_io_dina = {pipeline_1_out_addr,io_level}; // @[Cat.scala 30:58]
  assign buffer_io_wea = pipeline_1_m_axis_tvalid & pipeline_1_m_axis_tready; // @[BFS.scala 78:57]
  assign buffer_io_addrb = _buffer_io_addrb_T_8 | _buffer_io_addrb_T_7; // @[Mux.scala 27:72]
  assign buffer_io_clkb = clock; // @[BFS.scala 178:33]
  assign region_counter__addra = _region_counter_io_addra_T_1[9:0]; // @[BFS.scala 180:27]
  assign region_counter__clka = clock; // @[BFS.scala 54:41]
  assign region_counter__dina = _T_6 ? 9'h0 : region_counter_dina_0; // @[BFS.scala 182:32]
  assign region_counter__ena = 1'h1; // @[BFS.scala 55:25]
  assign region_counter__wea = _T_6 | _buffer_io_wea_T_2; // @[BFS.scala 181:31]
  assign region_counter__addrb = _region_counter_io_addrb_T_6[9:0]; // @[BFS.scala 183:27]
  assign region_counter__clkb = clock; // @[BFS.scala 53:41]
  assign region_counter__enb = 1'h1; // @[BFS.scala 56:25]
  assign region_counter_doutb_forward_aclk = clock; // @[BFS.scala 61:55]
  assign region_counter_doutb_forward_aresetn = ~reset; // @[BFS.scala 62:46]
  assign region_counter_doutb_forward_s_axis_tdata = {{7'd0}, region_counter_dina_0}; // @[BFS.scala 33:8]
  assign region_counter_doutb_forward_s_axis_tkeep = 2'h0;
  assign region_counter_doutb_forward_s_axis_tvalid = _region_counter_doutb_forward_io_s_axis_tvalid_T_2 &
    _buffer_io_wea_T_2; // @[BFS.scala 88:55]
  assign region_counter_doutb_forward_s_axis_tlast = 1'h0;
  assign region_counter_doutb_forward_m_axis_tready = wb_sm == 2'h0; // @[BFS.scala 116:58]
  assign pipeline_1_aclk = clock; // @[BFS.scala 71:37]
  assign pipeline_1_aresetn = ~reset; // @[BFS.scala 72:28]
  assign pipeline_1_s_axis_tdata = {{4'd0}, _pipeline_1_io_s_axis_tdata_T_1}; // @[Cat.scala 30:58]
  assign pipeline_1_s_axis_tkeep = 4'h0;
  assign pipeline_1_s_axis_tvalid = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 73:51]
  assign pipeline_1_s_axis_tlast = 1'h0;
  assign pipeline_1_m_axis_tready = wb_sm == 2'h0; // @[BFS.scala 115:40]
  assign aw_buffer_din = aw_buffer_reg_slice_m_axis_tdata + level_base_addr_reg; // @[BFS.scala 195:59]
  assign aw_buffer_wr_en = aw_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 194:22]
  assign aw_buffer_rd_en = io_axi_ddr_aw_ready; // @[BFS.scala 204:22]
  assign aw_buffer_clk = clock; // @[BFS.scala 192:35]
  assign aw_buffer_srst = reset; // @[BFS.scala 193:36]
  assign w_buffer_din = w_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 212:19]
  assign w_buffer_wr_en = w_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 211:21]
  assign w_buffer_rd_en = io_axi_ddr_w_ready; // @[BFS.scala 218:21]
  assign w_buffer_clk = clock; // @[BFS.scala 209:34]
  assign w_buffer_srst = reset; // @[BFS.scala 210:35]
  assign w_buffer_reg_slice_aclk = clock; // @[BFS.scala 110:45]
  assign w_buffer_reg_slice_aresetn = ~reset; // @[BFS.scala 111:36]
  assign w_buffer_reg_slice_s_axis_tdata = {{30'd0}, buffer_io_doutb[33:0]}; // @[BFS.scala 206:56]
  assign w_buffer_reg_slice_s_axis_tkeep = 8'h0;
  assign w_buffer_reg_slice_s_axis_tvalid = _T_6 & _T_7; // @[BFS.scala 207:64]
  assign w_buffer_reg_slice_s_axis_tlast = 1'h0;
  assign w_buffer_reg_slice_m_axis_tready = ~w_buffer_full; // @[util.scala 219:13]
  assign aw_buffer_reg_slice_aclk = clock; // @[BFS.scala 113:46]
  assign aw_buffer_reg_slice_aresetn = ~reset; // @[BFS.scala 114:37]
  assign aw_buffer_reg_slice_s_axis_tdata = {{38'd0}, _aw_buffer_reg_slice_io_s_axis_tdata_T_2}; // @[BFS.scala 45:53]
  assign aw_buffer_reg_slice_s_axis_tkeep = 8'h0;
  assign aw_buffer_reg_slice_s_axis_tvalid = _T_6 & _T_9; // @[BFS.scala 190:65]
  assign aw_buffer_reg_slice_s_axis_tlast = 1'h0;
  assign aw_buffer_reg_slice_m_axis_tready = ~aw_buffer_full; // @[util.scala 219:13]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 100:22]
      wb_sm <= 2'h0; // @[BFS.scala 100:22]
    end else if (flush_start) begin // @[BFS.scala 134:20]
      wb_sm <= 2'h3; // @[BFS.scala 135:11]
    end else if (_T) begin // @[BFS.scala 136:38]
      if (region_counter_doutb == 9'h0) begin // @[BFS.scala 137:39]
        wb_sm <= 2'h2; // @[BFS.scala 138:13]
      end else begin
        wb_sm <= 2'h1; // @[BFS.scala 140:13]
      end
    end else if (wb_start) begin // @[BFS.scala 142:23]
      wb_sm <= 2'h1; // @[BFS.scala 143:11]
    end else begin
      wb_sm <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 101:22]
      count <= 8'h0; // @[BFS.scala 101:22]
    end else if (_flush_start_T | _T_1) begin // @[BFS.scala 163:53]
      count <= 8'h1; // @[BFS.scala 164:11]
    end else if (_T_10) begin // @[BFS.scala 166:50]
      count <= _count_T_1; // @[BFS.scala 167:11]
    end
    if (reset) begin // @[BFS.scala 104:31]
      wb_block_index <= 10'h0; // @[BFS.scala 104:31]
    end else begin
      wb_block_index <= _GEN_4[9:0];
    end
    if (reset) begin // @[BFS.scala 106:23]
      size_b <= 8'h0; // @[BFS.scala 106:23]
    end else begin
      size_b <= _GEN_1[7:0];
    end
    if (reset) begin // @[BFS.scala 107:36]
      level_base_addr_reg <= 64'h0; // @[BFS.scala 107:36]
    end else begin
      level_base_addr_reg <= io_level_base_addr; // @[BFS.scala 117:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_sm = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  wb_block_index = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  size_b = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  level_base_addr_reg = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WB_engine_2(
  input          clock,
  input          reset,
  input          io_axi_ddr_aw_ready,
  output         io_axi_ddr_aw_valid,
  output [63:0]  io_axi_ddr_aw_bits_awaddr,
  output [5:0]   io_axi_ddr_aw_bits_awid,
  input          io_axi_ddr_w_ready,
  output         io_axi_ddr_w_valid,
  output [127:0] io_axi_ddr_w_bits_wdata,
  output [15:0]  io_axi_ddr_w_bits_wstrb,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [31:0]  io_xbar_in_bits_tdata,
  input  [63:0]  io_level_base_addr,
  input  [31:0]  io_level,
  output         io_end,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] buffer_io_addra; // @[BFS.scala 25:22]
  wire  buffer_io_clka; // @[BFS.scala 25:22]
  wire [47:0] buffer_io_dina; // @[BFS.scala 25:22]
  wire  buffer_io_wea; // @[BFS.scala 25:22]
  wire [15:0] buffer_io_addrb; // @[BFS.scala 25:22]
  wire  buffer_io_clkb; // @[BFS.scala 25:22]
  wire [47:0] buffer_io_doutb; // @[BFS.scala 25:22]
  wire [9:0] region_counter__addra; // @[BFS.scala 26:30]
  wire  region_counter__clka; // @[BFS.scala 26:30]
  wire [8:0] region_counter__dina; // @[BFS.scala 26:30]
  wire  region_counter__ena; // @[BFS.scala 26:30]
  wire  region_counter__wea; // @[BFS.scala 26:30]
  wire [9:0] region_counter__addrb; // @[BFS.scala 26:30]
  wire  region_counter__clkb; // @[BFS.scala 26:30]
  wire [8:0] region_counter__doutb; // @[BFS.scala 26:30]
  wire  region_counter__enb; // @[BFS.scala 26:30]
  wire  region_counter_doutb_forward_aclk; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_aresetn; // @[BFS.scala 60:44]
  wire [15:0] region_counter_doutb_forward_s_axis_tdata; // @[BFS.scala 60:44]
  wire [1:0] region_counter_doutb_forward_s_axis_tkeep; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tvalid; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tready; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tlast; // @[BFS.scala 60:44]
  wire [15:0] region_counter_doutb_forward_m_axis_tdata; // @[BFS.scala 60:44]
  wire [1:0] region_counter_doutb_forward_m_axis_tkeep; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tvalid; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tready; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tlast; // @[BFS.scala 60:44]
  wire  pipeline_1_aclk; // @[BFS.scala 64:26]
  wire  pipeline_1_aresetn; // @[BFS.scala 64:26]
  wire [31:0] pipeline_1_s_axis_tdata; // @[BFS.scala 64:26]
  wire [3:0] pipeline_1_s_axis_tkeep; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tvalid; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tready; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tlast; // @[BFS.scala 64:26]
  wire [31:0] pipeline_1_m_axis_tdata; // @[BFS.scala 64:26]
  wire [3:0] pipeline_1_m_axis_tkeep; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tvalid; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tready; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tlast; // @[BFS.scala 64:26]
  wire  aw_buffer_full; // @[BFS.scala 102:25]
  wire [63:0] aw_buffer_din; // @[BFS.scala 102:25]
  wire  aw_buffer_wr_en; // @[BFS.scala 102:25]
  wire  aw_buffer_empty; // @[BFS.scala 102:25]
  wire [63:0] aw_buffer_dout; // @[BFS.scala 102:25]
  wire  aw_buffer_rd_en; // @[BFS.scala 102:25]
  wire [5:0] aw_buffer_data_count; // @[BFS.scala 102:25]
  wire  aw_buffer_clk; // @[BFS.scala 102:25]
  wire  aw_buffer_srst; // @[BFS.scala 102:25]
  wire  aw_buffer_valid; // @[BFS.scala 102:25]
  wire  w_buffer_full; // @[BFS.scala 103:24]
  wire [63:0] w_buffer_din; // @[BFS.scala 103:24]
  wire  w_buffer_wr_en; // @[BFS.scala 103:24]
  wire  w_buffer_empty; // @[BFS.scala 103:24]
  wire [63:0] w_buffer_dout; // @[BFS.scala 103:24]
  wire  w_buffer_rd_en; // @[BFS.scala 103:24]
  wire [5:0] w_buffer_data_count; // @[BFS.scala 103:24]
  wire  w_buffer_clk; // @[BFS.scala 103:24]
  wire  w_buffer_srst; // @[BFS.scala 103:24]
  wire  w_buffer_valid; // @[BFS.scala 103:24]
  wire  w_buffer_reg_slice_aclk; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_aresetn; // @[BFS.scala 109:34]
  wire [63:0] w_buffer_reg_slice_s_axis_tdata; // @[BFS.scala 109:34]
  wire [7:0] w_buffer_reg_slice_s_axis_tkeep; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tvalid; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tready; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tlast; // @[BFS.scala 109:34]
  wire [63:0] w_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 109:34]
  wire [7:0] w_buffer_reg_slice_m_axis_tkeep; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tready; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tlast; // @[BFS.scala 109:34]
  wire  aw_buffer_reg_slice_aclk; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_aresetn; // @[BFS.scala 112:35]
  wire [63:0] aw_buffer_reg_slice_s_axis_tdata; // @[BFS.scala 112:35]
  wire [7:0] aw_buffer_reg_slice_s_axis_tkeep; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tvalid; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tready; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tlast; // @[BFS.scala 112:35]
  wire [63:0] aw_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 112:35]
  wire [7:0] aw_buffer_reg_slice_m_axis_tkeep; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tready; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tlast; // @[BFS.scala 112:35]
  wire [9:0] block_index = io_xbar_in_bits_tdata[23:14]; // @[BFS.scala 37:8]
  wire [15:0] pipeline_1_out_addr = pipeline_1_m_axis_tdata[27:12]; // @[BFS.scala 69:52]
  wire [11:0] pipeline_1_out_block_index = pipeline_1_m_axis_tdata[11:0]; // @[BFS.scala 70:59]
  wire  _pipeline_1_io_s_axis_tvalid_T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 73:51]
  wire [15:0] pipeline_1_io_s_axis_tdata_hi = {{4'd0}, io_xbar_in_bits_tdata[13:2]}; // @[BFS.scala 41:66 BFS.scala 41:66]
  wire [11:0] pipeline_1_io_s_axis_tdata_lo = {{2'd0}, block_index}; // @[BFS.scala 74:73 BFS.scala 74:73]
  wire [27:0] _pipeline_1_io_s_axis_tdata_T_1 = {pipeline_1_io_s_axis_tdata_hi,pipeline_1_io_s_axis_tdata_lo}; // @[Cat.scala 30:58]
  wire  _buffer_io_wea_T = pipeline_1_m_axis_tvalid; // @[BFS.scala 78:54]
  wire  _buffer_io_wea_T_2 = pipeline_1_m_axis_tvalid & pipeline_1_m_axis_tready; // @[BFS.scala 78:57]
  wire [15:0] _region_counter_doutb_T_1 = region_counter_doutb_forward_m_axis_tvalid ?
    region_counter_doutb_forward_m_axis_tdata : {{7'd0}, region_counter__doutb}; // @[BFS.scala 90:30]
  wire [8:0] region_counter_doutb = _region_counter_doutb_T_1[8:0]; // @[BFS.scala 63:34 BFS.scala 90:24]
  wire [5:0] buffer_io_addra_lo = region_counter_doutb[5:0]; // @[BFS.scala 29:35 BFS.scala 29:35]
  wire [17:0] _buffer_io_addra_T = {pipeline_1_out_block_index,buffer_io_addra_lo}; // @[Cat.scala 30:58]
  wire  _region_counter_dina_0_T = region_counter_doutb == 9'h3f; // @[BFS.scala 33:17]
  wire [8:0] _region_counter_dina_0_T_2 = region_counter_doutb + 9'h1; // @[BFS.scala 33:40]
  wire [8:0] region_counter_dina_0 = region_counter_doutb == 9'h3f ? 9'h0 : _region_counter_dina_0_T_2; // @[BFS.scala 33:8]
  wire  _region_counter_doutb_forward_io_s_axis_tvalid_T_1 = pipeline_1_out_block_index == pipeline_1_io_s_axis_tdata_lo
    ; // @[BFS.scala 88:28]
  wire  _region_counter_doutb_forward_io_s_axis_tvalid_T_2 = _pipeline_1_io_s_axis_tvalid_T &
    _region_counter_doutb_forward_io_s_axis_tvalid_T_1; // @[BFS.scala 87:89]
  reg [1:0] wb_sm; // @[BFS.scala 100:22]
  reg [7:0] count; // @[BFS.scala 101:22]
  reg [9:0] wb_block_index; // @[BFS.scala 104:31]
  wire  _flush_start_T = wb_sm == 2'h0; // @[BFS.scala 105:28]
  wire  flush_start = wb_sm == 2'h0 & io_flush; // @[BFS.scala 105:42]
  reg [7:0] size_b; // @[BFS.scala 106:23]
  reg [63:0] level_base_addr_reg; // @[BFS.scala 107:36]
  wire  wb_start = _buffer_io_wea_T & _region_counter_dina_0_T & _flush_start_T; // @[BFS.scala 108:89]
  wire  _T = wb_sm == 2'h3; // @[BFS.scala 121:20]
  wire [8:0] _GEN_0 = wb_sm == 2'h3 ? region_counter_doutb : {{1'd0}, size_b}; // @[BFS.scala 121:38 BFS.scala 122:12 BFS.scala 106:23]
  wire [8:0] _GEN_1 = wb_start ? 9'h40 : _GEN_0; // @[BFS.scala 119:17 BFS.scala 120:12]
  wire  _T_1 = wb_sm == 2'h2; // @[BFS.scala 129:20]
  wire  _T_2 = wb_block_index != 10'h3ff; // @[BFS.scala 129:55]
  wire [9:0] _wb_block_index_T_1 = wb_block_index + 10'h1; // @[BFS.scala 130:38]
  wire [9:0] _GEN_2 = wb_sm == 2'h2 & wb_block_index != 10'h3ff ? _wb_block_index_T_1 : wb_block_index; // @[BFS.scala 129:72 BFS.scala 130:20 BFS.scala 104:31]
  wire [9:0] _GEN_3 = flush_start ? 10'h0 : _GEN_2; // @[BFS.scala 127:26 BFS.scala 128:20]
  wire [11:0] _GEN_4 = wb_start ? pipeline_1_out_block_index : {{2'd0}, _GEN_3}; // @[BFS.scala 125:17 BFS.scala 126:20]
  wire  _T_6 = wb_sm == 2'h1; // @[BFS.scala 144:20]
  wire  _T_7 = aw_buffer_reg_slice_s_axis_tready; // @[BFS.scala 144:82]
  wire  _T_9 = w_buffer_reg_slice_s_axis_tready; // @[BFS.scala 145:47]
  wire  _T_10 = wb_sm == 2'h1 & aw_buffer_reg_slice_s_axis_tready & _T_9; // @[BFS.scala 144:85]
  wire [1:0] _GEN_6 = io_flush ? 2'h2 : 2'h0; // @[BFS.scala 147:21 BFS.scala 148:15 BFS.scala 150:15]
  wire [1:0] _GEN_7 = count == size_b ? _GEN_6 : 2'h1; // @[BFS.scala 146:27 BFS.scala 153:13]
  wire [1:0] _GEN_8 = _T_2 ? 2'h3 : 2'h0; // @[BFS.scala 156:42 BFS.scala 157:13 BFS.scala 159:13]
  wire [1:0] _GEN_9 = _T_1 ? _GEN_8 : wb_sm; // @[BFS.scala 155:38 BFS.scala 100:22]
  wire [1:0] _GEN_10 = _T_10 ? _GEN_7 : _GEN_9; // @[BFS.scala 145:51]
  wire [7:0] _count_T_1 = count + 8'h1; // @[BFS.scala 167:20]
  wire [15:0] _buffer_io_addrb_T = {block_index,6'h0}; // @[Cat.scala 30:58]
  wire [5:0] buffer_io_addrb_lo_2 = count[5:0]; // @[BFS.scala 29:35 BFS.scala 29:35]
  wire [15:0] _buffer_io_addrb_T_4 = {wb_block_index,buffer_io_addrb_lo_2}; // @[Cat.scala 30:58]
  wire [15:0] _buffer_io_addrb_T_5 = wb_start ? _buffer_io_addrb_T : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_6 = _T ? _buffer_io_addrb_T : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_7 = _T_6 ? _buffer_io_addrb_T_4 : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_8 = _buffer_io_addrb_T_5 | _buffer_io_addrb_T_6; // @[Mux.scala 27:72]
  wire [11:0] _region_counter_io_addra_T_1 = _T_6 ? {{2'd0}, wb_block_index} : pipeline_1_out_block_index; // @[BFS.scala 180:33]
  wire [11:0] _region_counter_io_addrb_T_4 = _T_6 ? pipeline_1_out_block_index : {{2'd0}, block_index}; // @[Mux.scala 98:16]
  wire [11:0] _region_counter_io_addrb_T_5 = flush_start ? 12'h0 : _region_counter_io_addrb_T_4; // @[Mux.scala 98:16]
  wire [11:0] _region_counter_io_addrb_T_6 = _T_1 ? {{2'd0}, _wb_block_index_T_1} : _region_counter_io_addrb_T_5; // @[Mux.scala 98:16]
  wire [11:0] aw_buffer_reg_slice_io_s_axis_tdata_lo = buffer_io_doutb[43:32]; // @[BFS.scala 45:43]
  wire [23:0] _aw_buffer_reg_slice_io_s_axis_tdata_T_1 = {wb_block_index,2'h2,aw_buffer_reg_slice_io_s_axis_tdata_lo}; // @[Cat.scala 30:58]
  wire [25:0] _aw_buffer_reg_slice_io_s_axis_tdata_T_2 = {_aw_buffer_reg_slice_io_s_axis_tdata_T_1, 2'h0}; // @[BFS.scala 45:53]
  wire [59:0] alignment_addr = aw_buffer_dout[63:4]; // @[BFS.scala 196:41]
  wire [4:0] io_axi_ddr_aw_bits_awid_lo = aw_buffer_data_count[4:0]; // @[BFS.scala 199:76 BFS.scala 199:76]
  wire [3:0] alignment_offset = {w_buffer_dout[33:32], 2'h0}; // @[BFS.scala 213:52]
  wire [7:0] _io_axi_ddr_w_bits_wdata_T_1 = 4'h8 * alignment_offset; // @[BFS.scala 214:84]
  wire [127:0] _io_axi_ddr_w_bits_wdata_WIRE = {{96'd0}, w_buffer_dout[31:0]}; // @[BFS.scala 214:62 BFS.scala 214:62]
  wire [382:0] _GEN_17 = {{255'd0}, _io_axi_ddr_w_bits_wdata_WIRE}; // @[BFS.scala 214:76]
  wire [382:0] _io_axi_ddr_w_bits_wdata_T_2 = _GEN_17 << _io_axi_ddr_w_bits_wdata_T_1; // @[BFS.scala 214:76]
  wire [30:0] _io_axi_ddr_w_bits_wstrb_T = 31'hf << alignment_offset; // @[BFS.scala 217:42]
  URAM_cluster buffer ( // @[BFS.scala 25:22]
    .io_addra(buffer_io_addra),
    .io_clka(buffer_io_clka),
    .io_dina(buffer_io_dina),
    .io_wea(buffer_io_wea),
    .io_addrb(buffer_io_addrb),
    .io_clkb(buffer_io_clkb),
    .io_doutb(buffer_io_doutb)
  );
  region_counter region_counter_ ( // @[BFS.scala 26:30]
    .addra(region_counter__addra),
    .clka(region_counter__clka),
    .dina(region_counter__dina),
    .ena(region_counter__ena),
    .wea(region_counter__wea),
    .addrb(region_counter__addrb),
    .clkb(region_counter__clkb),
    .doutb(region_counter__doutb),
    .enb(region_counter__enb)
  );
  region_counter_doutb_forward_reg_slice region_counter_doutb_forward ( // @[BFS.scala 60:44]
    .aclk(region_counter_doutb_forward_aclk),
    .aresetn(region_counter_doutb_forward_aresetn),
    .s_axis_tdata(region_counter_doutb_forward_s_axis_tdata),
    .s_axis_tkeep(region_counter_doutb_forward_s_axis_tkeep),
    .s_axis_tvalid(region_counter_doutb_forward_s_axis_tvalid),
    .s_axis_tready(region_counter_doutb_forward_s_axis_tready),
    .s_axis_tlast(region_counter_doutb_forward_s_axis_tlast),
    .m_axis_tdata(region_counter_doutb_forward_m_axis_tdata),
    .m_axis_tkeep(region_counter_doutb_forward_m_axis_tkeep),
    .m_axis_tvalid(region_counter_doutb_forward_m_axis_tvalid),
    .m_axis_tready(region_counter_doutb_forward_m_axis_tready),
    .m_axis_tlast(region_counter_doutb_forward_m_axis_tlast)
  );
  WB_engine_in_reg_slice pipeline_1 ( // @[BFS.scala 64:26]
    .aclk(pipeline_1_aclk),
    .aresetn(pipeline_1_aresetn),
    .s_axis_tdata(pipeline_1_s_axis_tdata),
    .s_axis_tkeep(pipeline_1_s_axis_tkeep),
    .s_axis_tvalid(pipeline_1_s_axis_tvalid),
    .s_axis_tready(pipeline_1_s_axis_tready),
    .s_axis_tlast(pipeline_1_s_axis_tlast),
    .m_axis_tdata(pipeline_1_m_axis_tdata),
    .m_axis_tkeep(pipeline_1_m_axis_tkeep),
    .m_axis_tvalid(pipeline_1_m_axis_tvalid),
    .m_axis_tready(pipeline_1_m_axis_tready),
    .m_axis_tlast(pipeline_1_m_axis_tlast)
  );
  addr_fifo aw_buffer ( // @[BFS.scala 102:25]
    .full(aw_buffer_full),
    .din(aw_buffer_din),
    .wr_en(aw_buffer_wr_en),
    .empty(aw_buffer_empty),
    .dout(aw_buffer_dout),
    .rd_en(aw_buffer_rd_en),
    .data_count(aw_buffer_data_count),
    .clk(aw_buffer_clk),
    .srst(aw_buffer_srst),
    .valid(aw_buffer_valid)
  );
  level_fifo w_buffer ( // @[BFS.scala 103:24]
    .full(w_buffer_full),
    .din(w_buffer_din),
    .wr_en(w_buffer_wr_en),
    .empty(w_buffer_empty),
    .dout(w_buffer_dout),
    .rd_en(w_buffer_rd_en),
    .data_count(w_buffer_data_count),
    .clk(w_buffer_clk),
    .srst(w_buffer_srst),
    .valid(w_buffer_valid)
  );
  w_buffer_reg_slice w_buffer_reg_slice ( // @[BFS.scala 109:34]
    .aclk(w_buffer_reg_slice_aclk),
    .aresetn(w_buffer_reg_slice_aresetn),
    .s_axis_tdata(w_buffer_reg_slice_s_axis_tdata),
    .s_axis_tkeep(w_buffer_reg_slice_s_axis_tkeep),
    .s_axis_tvalid(w_buffer_reg_slice_s_axis_tvalid),
    .s_axis_tready(w_buffer_reg_slice_s_axis_tready),
    .s_axis_tlast(w_buffer_reg_slice_s_axis_tlast),
    .m_axis_tdata(w_buffer_reg_slice_m_axis_tdata),
    .m_axis_tkeep(w_buffer_reg_slice_m_axis_tkeep),
    .m_axis_tvalid(w_buffer_reg_slice_m_axis_tvalid),
    .m_axis_tready(w_buffer_reg_slice_m_axis_tready),
    .m_axis_tlast(w_buffer_reg_slice_m_axis_tlast)
  );
  aw_buffer_reg_slice aw_buffer_reg_slice ( // @[BFS.scala 112:35]
    .aclk(aw_buffer_reg_slice_aclk),
    .aresetn(aw_buffer_reg_slice_aresetn),
    .s_axis_tdata(aw_buffer_reg_slice_s_axis_tdata),
    .s_axis_tkeep(aw_buffer_reg_slice_s_axis_tkeep),
    .s_axis_tvalid(aw_buffer_reg_slice_s_axis_tvalid),
    .s_axis_tready(aw_buffer_reg_slice_s_axis_tready),
    .s_axis_tlast(aw_buffer_reg_slice_s_axis_tlast),
    .m_axis_tdata(aw_buffer_reg_slice_m_axis_tdata),
    .m_axis_tkeep(aw_buffer_reg_slice_m_axis_tkeep),
    .m_axis_tvalid(aw_buffer_reg_slice_m_axis_tvalid),
    .m_axis_tready(aw_buffer_reg_slice_m_axis_tready),
    .m_axis_tlast(aw_buffer_reg_slice_m_axis_tlast)
  );
  assign io_axi_ddr_aw_valid = aw_buffer_valid; // @[BFS.scala 203:23]
  assign io_axi_ddr_aw_bits_awaddr = {alignment_addr,4'h0}; // @[Cat.scala 30:58]
  assign io_axi_ddr_aw_bits_awid = {1'h1,io_axi_ddr_aw_bits_awid_lo}; // @[Cat.scala 30:58]
  assign io_axi_ddr_w_valid = w_buffer_valid; // @[BFS.scala 216:22]
  assign io_axi_ddr_w_bits_wdata = _io_axi_ddr_w_bits_wdata_T_2[127:0]; // @[BFS.scala 214:27]
  assign io_axi_ddr_w_bits_wstrb = _io_axi_ddr_w_bits_wstrb_T[15:0]; // @[BFS.scala 217:27]
  assign io_xbar_in_ready = pipeline_1_s_axis_tready; // @[BFS.scala 75:20]
  assign io_end = _T_1 & wb_block_index == 10'h3ff; // @[BFS.scala 221:36]
  assign buffer_io_addra = _buffer_io_addra_T[15:0]; // @[BFS.scala 79:19]
  assign buffer_io_clka = clock; // @[BFS.scala 81:33]
  assign buffer_io_dina = {pipeline_1_out_addr,io_level}; // @[Cat.scala 30:58]
  assign buffer_io_wea = pipeline_1_m_axis_tvalid & pipeline_1_m_axis_tready; // @[BFS.scala 78:57]
  assign buffer_io_addrb = _buffer_io_addrb_T_8 | _buffer_io_addrb_T_7; // @[Mux.scala 27:72]
  assign buffer_io_clkb = clock; // @[BFS.scala 178:33]
  assign region_counter__addra = _region_counter_io_addra_T_1[9:0]; // @[BFS.scala 180:27]
  assign region_counter__clka = clock; // @[BFS.scala 54:41]
  assign region_counter__dina = _T_6 ? 9'h0 : region_counter_dina_0; // @[BFS.scala 182:32]
  assign region_counter__ena = 1'h1; // @[BFS.scala 55:25]
  assign region_counter__wea = _T_6 | _buffer_io_wea_T_2; // @[BFS.scala 181:31]
  assign region_counter__addrb = _region_counter_io_addrb_T_6[9:0]; // @[BFS.scala 183:27]
  assign region_counter__clkb = clock; // @[BFS.scala 53:41]
  assign region_counter__enb = 1'h1; // @[BFS.scala 56:25]
  assign region_counter_doutb_forward_aclk = clock; // @[BFS.scala 61:55]
  assign region_counter_doutb_forward_aresetn = ~reset; // @[BFS.scala 62:46]
  assign region_counter_doutb_forward_s_axis_tdata = {{7'd0}, region_counter_dina_0}; // @[BFS.scala 33:8]
  assign region_counter_doutb_forward_s_axis_tkeep = 2'h0;
  assign region_counter_doutb_forward_s_axis_tvalid = _region_counter_doutb_forward_io_s_axis_tvalid_T_2 &
    _buffer_io_wea_T_2; // @[BFS.scala 88:55]
  assign region_counter_doutb_forward_s_axis_tlast = 1'h0;
  assign region_counter_doutb_forward_m_axis_tready = wb_sm == 2'h0; // @[BFS.scala 116:58]
  assign pipeline_1_aclk = clock; // @[BFS.scala 71:37]
  assign pipeline_1_aresetn = ~reset; // @[BFS.scala 72:28]
  assign pipeline_1_s_axis_tdata = {{4'd0}, _pipeline_1_io_s_axis_tdata_T_1}; // @[Cat.scala 30:58]
  assign pipeline_1_s_axis_tkeep = 4'h0;
  assign pipeline_1_s_axis_tvalid = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 73:51]
  assign pipeline_1_s_axis_tlast = 1'h0;
  assign pipeline_1_m_axis_tready = wb_sm == 2'h0; // @[BFS.scala 115:40]
  assign aw_buffer_din = aw_buffer_reg_slice_m_axis_tdata + level_base_addr_reg; // @[BFS.scala 195:59]
  assign aw_buffer_wr_en = aw_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 194:22]
  assign aw_buffer_rd_en = io_axi_ddr_aw_ready; // @[BFS.scala 204:22]
  assign aw_buffer_clk = clock; // @[BFS.scala 192:35]
  assign aw_buffer_srst = reset; // @[BFS.scala 193:36]
  assign w_buffer_din = w_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 212:19]
  assign w_buffer_wr_en = w_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 211:21]
  assign w_buffer_rd_en = io_axi_ddr_w_ready; // @[BFS.scala 218:21]
  assign w_buffer_clk = clock; // @[BFS.scala 209:34]
  assign w_buffer_srst = reset; // @[BFS.scala 210:35]
  assign w_buffer_reg_slice_aclk = clock; // @[BFS.scala 110:45]
  assign w_buffer_reg_slice_aresetn = ~reset; // @[BFS.scala 111:36]
  assign w_buffer_reg_slice_s_axis_tdata = {{30'd0}, buffer_io_doutb[33:0]}; // @[BFS.scala 206:56]
  assign w_buffer_reg_slice_s_axis_tkeep = 8'h0;
  assign w_buffer_reg_slice_s_axis_tvalid = _T_6 & _T_7; // @[BFS.scala 207:64]
  assign w_buffer_reg_slice_s_axis_tlast = 1'h0;
  assign w_buffer_reg_slice_m_axis_tready = ~w_buffer_full; // @[util.scala 219:13]
  assign aw_buffer_reg_slice_aclk = clock; // @[BFS.scala 113:46]
  assign aw_buffer_reg_slice_aresetn = ~reset; // @[BFS.scala 114:37]
  assign aw_buffer_reg_slice_s_axis_tdata = {{38'd0}, _aw_buffer_reg_slice_io_s_axis_tdata_T_2}; // @[BFS.scala 45:53]
  assign aw_buffer_reg_slice_s_axis_tkeep = 8'h0;
  assign aw_buffer_reg_slice_s_axis_tvalid = _T_6 & _T_9; // @[BFS.scala 190:65]
  assign aw_buffer_reg_slice_s_axis_tlast = 1'h0;
  assign aw_buffer_reg_slice_m_axis_tready = ~aw_buffer_full; // @[util.scala 219:13]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 100:22]
      wb_sm <= 2'h0; // @[BFS.scala 100:22]
    end else if (flush_start) begin // @[BFS.scala 134:20]
      wb_sm <= 2'h3; // @[BFS.scala 135:11]
    end else if (_T) begin // @[BFS.scala 136:38]
      if (region_counter_doutb == 9'h0) begin // @[BFS.scala 137:39]
        wb_sm <= 2'h2; // @[BFS.scala 138:13]
      end else begin
        wb_sm <= 2'h1; // @[BFS.scala 140:13]
      end
    end else if (wb_start) begin // @[BFS.scala 142:23]
      wb_sm <= 2'h1; // @[BFS.scala 143:11]
    end else begin
      wb_sm <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 101:22]
      count <= 8'h0; // @[BFS.scala 101:22]
    end else if (_flush_start_T | _T_1) begin // @[BFS.scala 163:53]
      count <= 8'h1; // @[BFS.scala 164:11]
    end else if (_T_10) begin // @[BFS.scala 166:50]
      count <= _count_T_1; // @[BFS.scala 167:11]
    end
    if (reset) begin // @[BFS.scala 104:31]
      wb_block_index <= 10'h0; // @[BFS.scala 104:31]
    end else begin
      wb_block_index <= _GEN_4[9:0];
    end
    if (reset) begin // @[BFS.scala 106:23]
      size_b <= 8'h0; // @[BFS.scala 106:23]
    end else begin
      size_b <= _GEN_1[7:0];
    end
    if (reset) begin // @[BFS.scala 107:36]
      level_base_addr_reg <= 64'h0; // @[BFS.scala 107:36]
    end else begin
      level_base_addr_reg <= io_level_base_addr; // @[BFS.scala 117:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_sm = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  wb_block_index = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  size_b = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  level_base_addr_reg = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WB_engine_3(
  input          clock,
  input          reset,
  input          io_axi_ddr_aw_ready,
  output         io_axi_ddr_aw_valid,
  output [63:0]  io_axi_ddr_aw_bits_awaddr,
  output [5:0]   io_axi_ddr_aw_bits_awid,
  input          io_axi_ddr_w_ready,
  output         io_axi_ddr_w_valid,
  output [127:0] io_axi_ddr_w_bits_wdata,
  output [15:0]  io_axi_ddr_w_bits_wstrb,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [31:0]  io_xbar_in_bits_tdata,
  input  [63:0]  io_level_base_addr,
  input  [31:0]  io_level,
  output         io_end,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] buffer_io_addra; // @[BFS.scala 25:22]
  wire  buffer_io_clka; // @[BFS.scala 25:22]
  wire [47:0] buffer_io_dina; // @[BFS.scala 25:22]
  wire  buffer_io_wea; // @[BFS.scala 25:22]
  wire [15:0] buffer_io_addrb; // @[BFS.scala 25:22]
  wire  buffer_io_clkb; // @[BFS.scala 25:22]
  wire [47:0] buffer_io_doutb; // @[BFS.scala 25:22]
  wire [9:0] region_counter__addra; // @[BFS.scala 26:30]
  wire  region_counter__clka; // @[BFS.scala 26:30]
  wire [8:0] region_counter__dina; // @[BFS.scala 26:30]
  wire  region_counter__ena; // @[BFS.scala 26:30]
  wire  region_counter__wea; // @[BFS.scala 26:30]
  wire [9:0] region_counter__addrb; // @[BFS.scala 26:30]
  wire  region_counter__clkb; // @[BFS.scala 26:30]
  wire [8:0] region_counter__doutb; // @[BFS.scala 26:30]
  wire  region_counter__enb; // @[BFS.scala 26:30]
  wire  region_counter_doutb_forward_aclk; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_aresetn; // @[BFS.scala 60:44]
  wire [15:0] region_counter_doutb_forward_s_axis_tdata; // @[BFS.scala 60:44]
  wire [1:0] region_counter_doutb_forward_s_axis_tkeep; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tvalid; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tready; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_s_axis_tlast; // @[BFS.scala 60:44]
  wire [15:0] region_counter_doutb_forward_m_axis_tdata; // @[BFS.scala 60:44]
  wire [1:0] region_counter_doutb_forward_m_axis_tkeep; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tvalid; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tready; // @[BFS.scala 60:44]
  wire  region_counter_doutb_forward_m_axis_tlast; // @[BFS.scala 60:44]
  wire  pipeline_1_aclk; // @[BFS.scala 64:26]
  wire  pipeline_1_aresetn; // @[BFS.scala 64:26]
  wire [31:0] pipeline_1_s_axis_tdata; // @[BFS.scala 64:26]
  wire [3:0] pipeline_1_s_axis_tkeep; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tvalid; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tready; // @[BFS.scala 64:26]
  wire  pipeline_1_s_axis_tlast; // @[BFS.scala 64:26]
  wire [31:0] pipeline_1_m_axis_tdata; // @[BFS.scala 64:26]
  wire [3:0] pipeline_1_m_axis_tkeep; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tvalid; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tready; // @[BFS.scala 64:26]
  wire  pipeline_1_m_axis_tlast; // @[BFS.scala 64:26]
  wire  aw_buffer_full; // @[BFS.scala 102:25]
  wire [63:0] aw_buffer_din; // @[BFS.scala 102:25]
  wire  aw_buffer_wr_en; // @[BFS.scala 102:25]
  wire  aw_buffer_empty; // @[BFS.scala 102:25]
  wire [63:0] aw_buffer_dout; // @[BFS.scala 102:25]
  wire  aw_buffer_rd_en; // @[BFS.scala 102:25]
  wire [5:0] aw_buffer_data_count; // @[BFS.scala 102:25]
  wire  aw_buffer_clk; // @[BFS.scala 102:25]
  wire  aw_buffer_srst; // @[BFS.scala 102:25]
  wire  aw_buffer_valid; // @[BFS.scala 102:25]
  wire  w_buffer_full; // @[BFS.scala 103:24]
  wire [63:0] w_buffer_din; // @[BFS.scala 103:24]
  wire  w_buffer_wr_en; // @[BFS.scala 103:24]
  wire  w_buffer_empty; // @[BFS.scala 103:24]
  wire [63:0] w_buffer_dout; // @[BFS.scala 103:24]
  wire  w_buffer_rd_en; // @[BFS.scala 103:24]
  wire [5:0] w_buffer_data_count; // @[BFS.scala 103:24]
  wire  w_buffer_clk; // @[BFS.scala 103:24]
  wire  w_buffer_srst; // @[BFS.scala 103:24]
  wire  w_buffer_valid; // @[BFS.scala 103:24]
  wire  w_buffer_reg_slice_aclk; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_aresetn; // @[BFS.scala 109:34]
  wire [63:0] w_buffer_reg_slice_s_axis_tdata; // @[BFS.scala 109:34]
  wire [7:0] w_buffer_reg_slice_s_axis_tkeep; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tvalid; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tready; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_s_axis_tlast; // @[BFS.scala 109:34]
  wire [63:0] w_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 109:34]
  wire [7:0] w_buffer_reg_slice_m_axis_tkeep; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tready; // @[BFS.scala 109:34]
  wire  w_buffer_reg_slice_m_axis_tlast; // @[BFS.scala 109:34]
  wire  aw_buffer_reg_slice_aclk; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_aresetn; // @[BFS.scala 112:35]
  wire [63:0] aw_buffer_reg_slice_s_axis_tdata; // @[BFS.scala 112:35]
  wire [7:0] aw_buffer_reg_slice_s_axis_tkeep; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tvalid; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tready; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_s_axis_tlast; // @[BFS.scala 112:35]
  wire [63:0] aw_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 112:35]
  wire [7:0] aw_buffer_reg_slice_m_axis_tkeep; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tready; // @[BFS.scala 112:35]
  wire  aw_buffer_reg_slice_m_axis_tlast; // @[BFS.scala 112:35]
  wire [9:0] block_index = io_xbar_in_bits_tdata[23:14]; // @[BFS.scala 37:8]
  wire [15:0] pipeline_1_out_addr = pipeline_1_m_axis_tdata[27:12]; // @[BFS.scala 69:52]
  wire [11:0] pipeline_1_out_block_index = pipeline_1_m_axis_tdata[11:0]; // @[BFS.scala 70:59]
  wire  _pipeline_1_io_s_axis_tvalid_T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 73:51]
  wire [15:0] pipeline_1_io_s_axis_tdata_hi = {{4'd0}, io_xbar_in_bits_tdata[13:2]}; // @[BFS.scala 41:66 BFS.scala 41:66]
  wire [11:0] pipeline_1_io_s_axis_tdata_lo = {{2'd0}, block_index}; // @[BFS.scala 74:73 BFS.scala 74:73]
  wire [27:0] _pipeline_1_io_s_axis_tdata_T_1 = {pipeline_1_io_s_axis_tdata_hi,pipeline_1_io_s_axis_tdata_lo}; // @[Cat.scala 30:58]
  wire  _buffer_io_wea_T = pipeline_1_m_axis_tvalid; // @[BFS.scala 78:54]
  wire  _buffer_io_wea_T_2 = pipeline_1_m_axis_tvalid & pipeline_1_m_axis_tready; // @[BFS.scala 78:57]
  wire [15:0] _region_counter_doutb_T_1 = region_counter_doutb_forward_m_axis_tvalid ?
    region_counter_doutb_forward_m_axis_tdata : {{7'd0}, region_counter__doutb}; // @[BFS.scala 90:30]
  wire [8:0] region_counter_doutb = _region_counter_doutb_T_1[8:0]; // @[BFS.scala 63:34 BFS.scala 90:24]
  wire [5:0] buffer_io_addra_lo = region_counter_doutb[5:0]; // @[BFS.scala 29:35 BFS.scala 29:35]
  wire [17:0] _buffer_io_addra_T = {pipeline_1_out_block_index,buffer_io_addra_lo}; // @[Cat.scala 30:58]
  wire  _region_counter_dina_0_T = region_counter_doutb == 9'h3f; // @[BFS.scala 33:17]
  wire [8:0] _region_counter_dina_0_T_2 = region_counter_doutb + 9'h1; // @[BFS.scala 33:40]
  wire [8:0] region_counter_dina_0 = region_counter_doutb == 9'h3f ? 9'h0 : _region_counter_dina_0_T_2; // @[BFS.scala 33:8]
  wire  _region_counter_doutb_forward_io_s_axis_tvalid_T_1 = pipeline_1_out_block_index == pipeline_1_io_s_axis_tdata_lo
    ; // @[BFS.scala 88:28]
  wire  _region_counter_doutb_forward_io_s_axis_tvalid_T_2 = _pipeline_1_io_s_axis_tvalid_T &
    _region_counter_doutb_forward_io_s_axis_tvalid_T_1; // @[BFS.scala 87:89]
  reg [1:0] wb_sm; // @[BFS.scala 100:22]
  reg [7:0] count; // @[BFS.scala 101:22]
  reg [9:0] wb_block_index; // @[BFS.scala 104:31]
  wire  _flush_start_T = wb_sm == 2'h0; // @[BFS.scala 105:28]
  wire  flush_start = wb_sm == 2'h0 & io_flush; // @[BFS.scala 105:42]
  reg [7:0] size_b; // @[BFS.scala 106:23]
  reg [63:0] level_base_addr_reg; // @[BFS.scala 107:36]
  wire  wb_start = _buffer_io_wea_T & _region_counter_dina_0_T & _flush_start_T; // @[BFS.scala 108:89]
  wire  _T = wb_sm == 2'h3; // @[BFS.scala 121:20]
  wire [8:0] _GEN_0 = wb_sm == 2'h3 ? region_counter_doutb : {{1'd0}, size_b}; // @[BFS.scala 121:38 BFS.scala 122:12 BFS.scala 106:23]
  wire [8:0] _GEN_1 = wb_start ? 9'h40 : _GEN_0; // @[BFS.scala 119:17 BFS.scala 120:12]
  wire  _T_1 = wb_sm == 2'h2; // @[BFS.scala 129:20]
  wire  _T_2 = wb_block_index != 10'h3ff; // @[BFS.scala 129:55]
  wire [9:0] _wb_block_index_T_1 = wb_block_index + 10'h1; // @[BFS.scala 130:38]
  wire [9:0] _GEN_2 = wb_sm == 2'h2 & wb_block_index != 10'h3ff ? _wb_block_index_T_1 : wb_block_index; // @[BFS.scala 129:72 BFS.scala 130:20 BFS.scala 104:31]
  wire [9:0] _GEN_3 = flush_start ? 10'h0 : _GEN_2; // @[BFS.scala 127:26 BFS.scala 128:20]
  wire [11:0] _GEN_4 = wb_start ? pipeline_1_out_block_index : {{2'd0}, _GEN_3}; // @[BFS.scala 125:17 BFS.scala 126:20]
  wire  _T_6 = wb_sm == 2'h1; // @[BFS.scala 144:20]
  wire  _T_7 = aw_buffer_reg_slice_s_axis_tready; // @[BFS.scala 144:82]
  wire  _T_9 = w_buffer_reg_slice_s_axis_tready; // @[BFS.scala 145:47]
  wire  _T_10 = wb_sm == 2'h1 & aw_buffer_reg_slice_s_axis_tready & _T_9; // @[BFS.scala 144:85]
  wire [1:0] _GEN_6 = io_flush ? 2'h2 : 2'h0; // @[BFS.scala 147:21 BFS.scala 148:15 BFS.scala 150:15]
  wire [1:0] _GEN_7 = count == size_b ? _GEN_6 : 2'h1; // @[BFS.scala 146:27 BFS.scala 153:13]
  wire [1:0] _GEN_8 = _T_2 ? 2'h3 : 2'h0; // @[BFS.scala 156:42 BFS.scala 157:13 BFS.scala 159:13]
  wire [1:0] _GEN_9 = _T_1 ? _GEN_8 : wb_sm; // @[BFS.scala 155:38 BFS.scala 100:22]
  wire [1:0] _GEN_10 = _T_10 ? _GEN_7 : _GEN_9; // @[BFS.scala 145:51]
  wire [7:0] _count_T_1 = count + 8'h1; // @[BFS.scala 167:20]
  wire [15:0] _buffer_io_addrb_T = {block_index,6'h0}; // @[Cat.scala 30:58]
  wire [5:0] buffer_io_addrb_lo_2 = count[5:0]; // @[BFS.scala 29:35 BFS.scala 29:35]
  wire [15:0] _buffer_io_addrb_T_4 = {wb_block_index,buffer_io_addrb_lo_2}; // @[Cat.scala 30:58]
  wire [15:0] _buffer_io_addrb_T_5 = wb_start ? _buffer_io_addrb_T : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_6 = _T ? _buffer_io_addrb_T : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_7 = _T_6 ? _buffer_io_addrb_T_4 : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _buffer_io_addrb_T_8 = _buffer_io_addrb_T_5 | _buffer_io_addrb_T_6; // @[Mux.scala 27:72]
  wire [11:0] _region_counter_io_addra_T_1 = _T_6 ? {{2'd0}, wb_block_index} : pipeline_1_out_block_index; // @[BFS.scala 180:33]
  wire [11:0] _region_counter_io_addrb_T_4 = _T_6 ? pipeline_1_out_block_index : {{2'd0}, block_index}; // @[Mux.scala 98:16]
  wire [11:0] _region_counter_io_addrb_T_5 = flush_start ? 12'h0 : _region_counter_io_addrb_T_4; // @[Mux.scala 98:16]
  wire [11:0] _region_counter_io_addrb_T_6 = _T_1 ? {{2'd0}, _wb_block_index_T_1} : _region_counter_io_addrb_T_5; // @[Mux.scala 98:16]
  wire [11:0] aw_buffer_reg_slice_io_s_axis_tdata_lo = buffer_io_doutb[43:32]; // @[BFS.scala 45:43]
  wire [23:0] _aw_buffer_reg_slice_io_s_axis_tdata_T_1 = {wb_block_index,2'h3,aw_buffer_reg_slice_io_s_axis_tdata_lo}; // @[Cat.scala 30:58]
  wire [25:0] _aw_buffer_reg_slice_io_s_axis_tdata_T_2 = {_aw_buffer_reg_slice_io_s_axis_tdata_T_1, 2'h0}; // @[BFS.scala 45:53]
  wire [59:0] alignment_addr = aw_buffer_dout[63:4]; // @[BFS.scala 196:41]
  wire [4:0] io_axi_ddr_aw_bits_awid_lo = aw_buffer_data_count[4:0]; // @[BFS.scala 199:76 BFS.scala 199:76]
  wire [3:0] alignment_offset = {w_buffer_dout[33:32], 2'h0}; // @[BFS.scala 213:52]
  wire [7:0] _io_axi_ddr_w_bits_wdata_T_1 = 4'h8 * alignment_offset; // @[BFS.scala 214:84]
  wire [127:0] _io_axi_ddr_w_bits_wdata_WIRE = {{96'd0}, w_buffer_dout[31:0]}; // @[BFS.scala 214:62 BFS.scala 214:62]
  wire [382:0] _GEN_17 = {{255'd0}, _io_axi_ddr_w_bits_wdata_WIRE}; // @[BFS.scala 214:76]
  wire [382:0] _io_axi_ddr_w_bits_wdata_T_2 = _GEN_17 << _io_axi_ddr_w_bits_wdata_T_1; // @[BFS.scala 214:76]
  wire [30:0] _io_axi_ddr_w_bits_wstrb_T = 31'hf << alignment_offset; // @[BFS.scala 217:42]
  URAM_cluster buffer ( // @[BFS.scala 25:22]
    .io_addra(buffer_io_addra),
    .io_clka(buffer_io_clka),
    .io_dina(buffer_io_dina),
    .io_wea(buffer_io_wea),
    .io_addrb(buffer_io_addrb),
    .io_clkb(buffer_io_clkb),
    .io_doutb(buffer_io_doutb)
  );
  region_counter region_counter_ ( // @[BFS.scala 26:30]
    .addra(region_counter__addra),
    .clka(region_counter__clka),
    .dina(region_counter__dina),
    .ena(region_counter__ena),
    .wea(region_counter__wea),
    .addrb(region_counter__addrb),
    .clkb(region_counter__clkb),
    .doutb(region_counter__doutb),
    .enb(region_counter__enb)
  );
  region_counter_doutb_forward_reg_slice region_counter_doutb_forward ( // @[BFS.scala 60:44]
    .aclk(region_counter_doutb_forward_aclk),
    .aresetn(region_counter_doutb_forward_aresetn),
    .s_axis_tdata(region_counter_doutb_forward_s_axis_tdata),
    .s_axis_tkeep(region_counter_doutb_forward_s_axis_tkeep),
    .s_axis_tvalid(region_counter_doutb_forward_s_axis_tvalid),
    .s_axis_tready(region_counter_doutb_forward_s_axis_tready),
    .s_axis_tlast(region_counter_doutb_forward_s_axis_tlast),
    .m_axis_tdata(region_counter_doutb_forward_m_axis_tdata),
    .m_axis_tkeep(region_counter_doutb_forward_m_axis_tkeep),
    .m_axis_tvalid(region_counter_doutb_forward_m_axis_tvalid),
    .m_axis_tready(region_counter_doutb_forward_m_axis_tready),
    .m_axis_tlast(region_counter_doutb_forward_m_axis_tlast)
  );
  WB_engine_in_reg_slice pipeline_1 ( // @[BFS.scala 64:26]
    .aclk(pipeline_1_aclk),
    .aresetn(pipeline_1_aresetn),
    .s_axis_tdata(pipeline_1_s_axis_tdata),
    .s_axis_tkeep(pipeline_1_s_axis_tkeep),
    .s_axis_tvalid(pipeline_1_s_axis_tvalid),
    .s_axis_tready(pipeline_1_s_axis_tready),
    .s_axis_tlast(pipeline_1_s_axis_tlast),
    .m_axis_tdata(pipeline_1_m_axis_tdata),
    .m_axis_tkeep(pipeline_1_m_axis_tkeep),
    .m_axis_tvalid(pipeline_1_m_axis_tvalid),
    .m_axis_tready(pipeline_1_m_axis_tready),
    .m_axis_tlast(pipeline_1_m_axis_tlast)
  );
  addr_fifo aw_buffer ( // @[BFS.scala 102:25]
    .full(aw_buffer_full),
    .din(aw_buffer_din),
    .wr_en(aw_buffer_wr_en),
    .empty(aw_buffer_empty),
    .dout(aw_buffer_dout),
    .rd_en(aw_buffer_rd_en),
    .data_count(aw_buffer_data_count),
    .clk(aw_buffer_clk),
    .srst(aw_buffer_srst),
    .valid(aw_buffer_valid)
  );
  level_fifo w_buffer ( // @[BFS.scala 103:24]
    .full(w_buffer_full),
    .din(w_buffer_din),
    .wr_en(w_buffer_wr_en),
    .empty(w_buffer_empty),
    .dout(w_buffer_dout),
    .rd_en(w_buffer_rd_en),
    .data_count(w_buffer_data_count),
    .clk(w_buffer_clk),
    .srst(w_buffer_srst),
    .valid(w_buffer_valid)
  );
  w_buffer_reg_slice w_buffer_reg_slice ( // @[BFS.scala 109:34]
    .aclk(w_buffer_reg_slice_aclk),
    .aresetn(w_buffer_reg_slice_aresetn),
    .s_axis_tdata(w_buffer_reg_slice_s_axis_tdata),
    .s_axis_tkeep(w_buffer_reg_slice_s_axis_tkeep),
    .s_axis_tvalid(w_buffer_reg_slice_s_axis_tvalid),
    .s_axis_tready(w_buffer_reg_slice_s_axis_tready),
    .s_axis_tlast(w_buffer_reg_slice_s_axis_tlast),
    .m_axis_tdata(w_buffer_reg_slice_m_axis_tdata),
    .m_axis_tkeep(w_buffer_reg_slice_m_axis_tkeep),
    .m_axis_tvalid(w_buffer_reg_slice_m_axis_tvalid),
    .m_axis_tready(w_buffer_reg_slice_m_axis_tready),
    .m_axis_tlast(w_buffer_reg_slice_m_axis_tlast)
  );
  aw_buffer_reg_slice aw_buffer_reg_slice ( // @[BFS.scala 112:35]
    .aclk(aw_buffer_reg_slice_aclk),
    .aresetn(aw_buffer_reg_slice_aresetn),
    .s_axis_tdata(aw_buffer_reg_slice_s_axis_tdata),
    .s_axis_tkeep(aw_buffer_reg_slice_s_axis_tkeep),
    .s_axis_tvalid(aw_buffer_reg_slice_s_axis_tvalid),
    .s_axis_tready(aw_buffer_reg_slice_s_axis_tready),
    .s_axis_tlast(aw_buffer_reg_slice_s_axis_tlast),
    .m_axis_tdata(aw_buffer_reg_slice_m_axis_tdata),
    .m_axis_tkeep(aw_buffer_reg_slice_m_axis_tkeep),
    .m_axis_tvalid(aw_buffer_reg_slice_m_axis_tvalid),
    .m_axis_tready(aw_buffer_reg_slice_m_axis_tready),
    .m_axis_tlast(aw_buffer_reg_slice_m_axis_tlast)
  );
  assign io_axi_ddr_aw_valid = aw_buffer_valid; // @[BFS.scala 203:23]
  assign io_axi_ddr_aw_bits_awaddr = {alignment_addr,4'h0}; // @[Cat.scala 30:58]
  assign io_axi_ddr_aw_bits_awid = {1'h1,io_axi_ddr_aw_bits_awid_lo}; // @[Cat.scala 30:58]
  assign io_axi_ddr_w_valid = w_buffer_valid; // @[BFS.scala 216:22]
  assign io_axi_ddr_w_bits_wdata = _io_axi_ddr_w_bits_wdata_T_2[127:0]; // @[BFS.scala 214:27]
  assign io_axi_ddr_w_bits_wstrb = _io_axi_ddr_w_bits_wstrb_T[15:0]; // @[BFS.scala 217:27]
  assign io_xbar_in_ready = pipeline_1_s_axis_tready; // @[BFS.scala 75:20]
  assign io_end = _T_1 & wb_block_index == 10'h3ff; // @[BFS.scala 221:36]
  assign buffer_io_addra = _buffer_io_addra_T[15:0]; // @[BFS.scala 79:19]
  assign buffer_io_clka = clock; // @[BFS.scala 81:33]
  assign buffer_io_dina = {pipeline_1_out_addr,io_level}; // @[Cat.scala 30:58]
  assign buffer_io_wea = pipeline_1_m_axis_tvalid & pipeline_1_m_axis_tready; // @[BFS.scala 78:57]
  assign buffer_io_addrb = _buffer_io_addrb_T_8 | _buffer_io_addrb_T_7; // @[Mux.scala 27:72]
  assign buffer_io_clkb = clock; // @[BFS.scala 178:33]
  assign region_counter__addra = _region_counter_io_addra_T_1[9:0]; // @[BFS.scala 180:27]
  assign region_counter__clka = clock; // @[BFS.scala 54:41]
  assign region_counter__dina = _T_6 ? 9'h0 : region_counter_dina_0; // @[BFS.scala 182:32]
  assign region_counter__ena = 1'h1; // @[BFS.scala 55:25]
  assign region_counter__wea = _T_6 | _buffer_io_wea_T_2; // @[BFS.scala 181:31]
  assign region_counter__addrb = _region_counter_io_addrb_T_6[9:0]; // @[BFS.scala 183:27]
  assign region_counter__clkb = clock; // @[BFS.scala 53:41]
  assign region_counter__enb = 1'h1; // @[BFS.scala 56:25]
  assign region_counter_doutb_forward_aclk = clock; // @[BFS.scala 61:55]
  assign region_counter_doutb_forward_aresetn = ~reset; // @[BFS.scala 62:46]
  assign region_counter_doutb_forward_s_axis_tdata = {{7'd0}, region_counter_dina_0}; // @[BFS.scala 33:8]
  assign region_counter_doutb_forward_s_axis_tkeep = 2'h0;
  assign region_counter_doutb_forward_s_axis_tvalid = _region_counter_doutb_forward_io_s_axis_tvalid_T_2 &
    _buffer_io_wea_T_2; // @[BFS.scala 88:55]
  assign region_counter_doutb_forward_s_axis_tlast = 1'h0;
  assign region_counter_doutb_forward_m_axis_tready = wb_sm == 2'h0; // @[BFS.scala 116:58]
  assign pipeline_1_aclk = clock; // @[BFS.scala 71:37]
  assign pipeline_1_aresetn = ~reset; // @[BFS.scala 72:28]
  assign pipeline_1_s_axis_tdata = {{4'd0}, _pipeline_1_io_s_axis_tdata_T_1}; // @[Cat.scala 30:58]
  assign pipeline_1_s_axis_tkeep = 4'h0;
  assign pipeline_1_s_axis_tvalid = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 73:51]
  assign pipeline_1_s_axis_tlast = 1'h0;
  assign pipeline_1_m_axis_tready = wb_sm == 2'h0; // @[BFS.scala 115:40]
  assign aw_buffer_din = aw_buffer_reg_slice_m_axis_tdata + level_base_addr_reg; // @[BFS.scala 195:59]
  assign aw_buffer_wr_en = aw_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 194:22]
  assign aw_buffer_rd_en = io_axi_ddr_aw_ready; // @[BFS.scala 204:22]
  assign aw_buffer_clk = clock; // @[BFS.scala 192:35]
  assign aw_buffer_srst = reset; // @[BFS.scala 193:36]
  assign w_buffer_din = w_buffer_reg_slice_m_axis_tdata; // @[BFS.scala 212:19]
  assign w_buffer_wr_en = w_buffer_reg_slice_m_axis_tvalid; // @[BFS.scala 211:21]
  assign w_buffer_rd_en = io_axi_ddr_w_ready; // @[BFS.scala 218:21]
  assign w_buffer_clk = clock; // @[BFS.scala 209:34]
  assign w_buffer_srst = reset; // @[BFS.scala 210:35]
  assign w_buffer_reg_slice_aclk = clock; // @[BFS.scala 110:45]
  assign w_buffer_reg_slice_aresetn = ~reset; // @[BFS.scala 111:36]
  assign w_buffer_reg_slice_s_axis_tdata = {{30'd0}, buffer_io_doutb[33:0]}; // @[BFS.scala 206:56]
  assign w_buffer_reg_slice_s_axis_tkeep = 8'h0;
  assign w_buffer_reg_slice_s_axis_tvalid = _T_6 & _T_7; // @[BFS.scala 207:64]
  assign w_buffer_reg_slice_s_axis_tlast = 1'h0;
  assign w_buffer_reg_slice_m_axis_tready = ~w_buffer_full; // @[util.scala 219:13]
  assign aw_buffer_reg_slice_aclk = clock; // @[BFS.scala 113:46]
  assign aw_buffer_reg_slice_aresetn = ~reset; // @[BFS.scala 114:37]
  assign aw_buffer_reg_slice_s_axis_tdata = {{38'd0}, _aw_buffer_reg_slice_io_s_axis_tdata_T_2}; // @[BFS.scala 45:53]
  assign aw_buffer_reg_slice_s_axis_tkeep = 8'h0;
  assign aw_buffer_reg_slice_s_axis_tvalid = _T_6 & _T_9; // @[BFS.scala 190:65]
  assign aw_buffer_reg_slice_s_axis_tlast = 1'h0;
  assign aw_buffer_reg_slice_m_axis_tready = ~aw_buffer_full; // @[util.scala 219:13]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 100:22]
      wb_sm <= 2'h0; // @[BFS.scala 100:22]
    end else if (flush_start) begin // @[BFS.scala 134:20]
      wb_sm <= 2'h3; // @[BFS.scala 135:11]
    end else if (_T) begin // @[BFS.scala 136:38]
      if (region_counter_doutb == 9'h0) begin // @[BFS.scala 137:39]
        wb_sm <= 2'h2; // @[BFS.scala 138:13]
      end else begin
        wb_sm <= 2'h1; // @[BFS.scala 140:13]
      end
    end else if (wb_start) begin // @[BFS.scala 142:23]
      wb_sm <= 2'h1; // @[BFS.scala 143:11]
    end else begin
      wb_sm <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 101:22]
      count <= 8'h0; // @[BFS.scala 101:22]
    end else if (_flush_start_T | _T_1) begin // @[BFS.scala 163:53]
      count <= 8'h1; // @[BFS.scala 164:11]
    end else if (_T_10) begin // @[BFS.scala 166:50]
      count <= _count_T_1; // @[BFS.scala 167:11]
    end
    if (reset) begin // @[BFS.scala 104:31]
      wb_block_index <= 10'h0; // @[BFS.scala 104:31]
    end else begin
      wb_block_index <= _GEN_4[9:0];
    end
    if (reset) begin // @[BFS.scala 106:23]
      size_b <= 8'h0; // @[BFS.scala 106:23]
    end else begin
      size_b <= _GEN_1[7:0];
    end
    if (reset) begin // @[BFS.scala 107:36]
      level_base_addr_reg <= 64'h0; // @[BFS.scala 107:36]
    end else begin
      level_base_addr_reg <= io_level_base_addr; // @[BFS.scala 117:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_sm = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  wb_block_index = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  size_b = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  level_base_addr_reg = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Apply(
  input          clock,
  input          reset,
  input          io_axi_0_ddr_aw_ready,
  output         io_axi_0_ddr_aw_valid,
  output [63:0]  io_axi_0_ddr_aw_bits_awaddr,
  output [5:0]   io_axi_0_ddr_aw_bits_awid,
  input          io_axi_0_ddr_w_ready,
  output         io_axi_0_ddr_w_valid,
  output [127:0] io_axi_0_ddr_w_bits_wdata,
  output [15:0]  io_axi_0_ddr_w_bits_wstrb,
  input          io_axi_1_ddr_aw_ready,
  output         io_axi_1_ddr_aw_valid,
  output [63:0]  io_axi_1_ddr_aw_bits_awaddr,
  output [5:0]   io_axi_1_ddr_aw_bits_awid,
  input          io_axi_1_ddr_w_ready,
  output         io_axi_1_ddr_w_valid,
  output [127:0] io_axi_1_ddr_w_bits_wdata,
  output [15:0]  io_axi_1_ddr_w_bits_wstrb,
  input          io_axi_2_ddr_aw_ready,
  output         io_axi_2_ddr_aw_valid,
  output [63:0]  io_axi_2_ddr_aw_bits_awaddr,
  output [5:0]   io_axi_2_ddr_aw_bits_awid,
  input          io_axi_2_ddr_w_ready,
  output         io_axi_2_ddr_w_valid,
  output [127:0] io_axi_2_ddr_w_bits_wdata,
  output [15:0]  io_axi_2_ddr_w_bits_wstrb,
  input          io_axi_3_ddr_aw_ready,
  output         io_axi_3_ddr_aw_valid,
  output [63:0]  io_axi_3_ddr_aw_bits_awaddr,
  output [5:0]   io_axi_3_ddr_aw_bits_awid,
  input          io_axi_3_ddr_w_ready,
  output         io_axi_3_ddr_w_valid,
  output [127:0] io_axi_3_ddr_w_bits_wdata,
  output [15:0]  io_axi_3_ddr_w_bits_wstrb,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [511:0] io_gather_in_bits_tdata,
  input  [63:0]  io_gather_in_bits_tkeep,
  input          io_gather_in_bits_tlast,
  input  [31:0]  io_level,
  input  [63:0]  io_level_base_addr,
  output         io_end,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  apply_in_aclk; // @[BFS.scala 251:24]
  wire  apply_in_aresetn; // @[BFS.scala 251:24]
  wire [511:0] apply_in_s_axis_tdata; // @[BFS.scala 251:24]
  wire [63:0] apply_in_s_axis_tkeep; // @[BFS.scala 251:24]
  wire  apply_in_s_axis_tvalid; // @[BFS.scala 251:24]
  wire  apply_in_s_axis_tready; // @[BFS.scala 251:24]
  wire  apply_in_s_axis_tlast; // @[BFS.scala 251:24]
  wire [511:0] apply_in_m_axis_tdata; // @[BFS.scala 251:24]
  wire [63:0] apply_in_m_axis_tkeep; // @[BFS.scala 251:24]
  wire  apply_in_m_axis_tvalid; // @[BFS.scala 251:24]
  wire  apply_in_m_axis_tready; // @[BFS.scala 251:24]
  wire  apply_in_m_axis_tlast; // @[BFS.scala 251:24]
  wire  broadcaster_aclk; // @[BFS.scala 258:27]
  wire  broadcaster_aresetn; // @[BFS.scala 258:27]
  wire [511:0] broadcaster_s_axis_tdata; // @[BFS.scala 258:27]
  wire [63:0] broadcaster_s_axis_tkeep; // @[BFS.scala 258:27]
  wire  broadcaster_s_axis_tvalid; // @[BFS.scala 258:27]
  wire  broadcaster_s_axis_tready; // @[BFS.scala 258:27]
  wire  broadcaster_s_axis_tlast; // @[BFS.scala 258:27]
  wire  broadcaster_s_axis_tid; // @[BFS.scala 258:27]
  wire [2047:0] broadcaster_m_axis_tdata; // @[BFS.scala 258:27]
  wire [255:0] broadcaster_m_axis_tkeep; // @[BFS.scala 258:27]
  wire [3:0] broadcaster_m_axis_tvalid; // @[BFS.scala 258:27]
  wire [3:0] broadcaster_m_axis_tready; // @[BFS.scala 258:27]
  wire [3:0] broadcaster_m_axis_tlast; // @[BFS.scala 258:27]
  wire [3:0] broadcaster_m_axis_tid; // @[BFS.scala 258:27]
  wire  apply_selecter_0_clock; // @[BFS.scala 268:11]
  wire  apply_selecter_0_reset; // @[BFS.scala 268:11]
  wire  apply_selecter_0_io_xbar_in_ready; // @[BFS.scala 268:11]
  wire  apply_selecter_0_io_xbar_in_valid; // @[BFS.scala 268:11]
  wire [511:0] apply_selecter_0_io_xbar_in_bits_tdata; // @[BFS.scala 268:11]
  wire [15:0] apply_selecter_0_io_xbar_in_bits_tkeep; // @[BFS.scala 268:11]
  wire  apply_selecter_0_io_xbar_in_bits_tlast; // @[BFS.scala 268:11]
  wire  apply_selecter_0_io_ddr_out_ready; // @[BFS.scala 268:11]
  wire  apply_selecter_0_io_ddr_out_valid; // @[BFS.scala 268:11]
  wire [31:0] apply_selecter_0_io_ddr_out_bits_tdata; // @[BFS.scala 268:11]
  wire  apply_selecter_1_clock; // @[BFS.scala 268:11]
  wire  apply_selecter_1_reset; // @[BFS.scala 268:11]
  wire  apply_selecter_1_io_xbar_in_ready; // @[BFS.scala 268:11]
  wire  apply_selecter_1_io_xbar_in_valid; // @[BFS.scala 268:11]
  wire [511:0] apply_selecter_1_io_xbar_in_bits_tdata; // @[BFS.scala 268:11]
  wire [15:0] apply_selecter_1_io_xbar_in_bits_tkeep; // @[BFS.scala 268:11]
  wire  apply_selecter_1_io_xbar_in_bits_tlast; // @[BFS.scala 268:11]
  wire  apply_selecter_1_io_ddr_out_ready; // @[BFS.scala 268:11]
  wire  apply_selecter_1_io_ddr_out_valid; // @[BFS.scala 268:11]
  wire [31:0] apply_selecter_1_io_ddr_out_bits_tdata; // @[BFS.scala 268:11]
  wire  apply_selecter_2_clock; // @[BFS.scala 268:11]
  wire  apply_selecter_2_reset; // @[BFS.scala 268:11]
  wire  apply_selecter_2_io_xbar_in_ready; // @[BFS.scala 268:11]
  wire  apply_selecter_2_io_xbar_in_valid; // @[BFS.scala 268:11]
  wire [511:0] apply_selecter_2_io_xbar_in_bits_tdata; // @[BFS.scala 268:11]
  wire [15:0] apply_selecter_2_io_xbar_in_bits_tkeep; // @[BFS.scala 268:11]
  wire  apply_selecter_2_io_xbar_in_bits_tlast; // @[BFS.scala 268:11]
  wire  apply_selecter_2_io_ddr_out_ready; // @[BFS.scala 268:11]
  wire  apply_selecter_2_io_ddr_out_valid; // @[BFS.scala 268:11]
  wire [31:0] apply_selecter_2_io_ddr_out_bits_tdata; // @[BFS.scala 268:11]
  wire  apply_selecter_3_clock; // @[BFS.scala 268:11]
  wire  apply_selecter_3_reset; // @[BFS.scala 268:11]
  wire  apply_selecter_3_io_xbar_in_ready; // @[BFS.scala 268:11]
  wire  apply_selecter_3_io_xbar_in_valid; // @[BFS.scala 268:11]
  wire [511:0] apply_selecter_3_io_xbar_in_bits_tdata; // @[BFS.scala 268:11]
  wire [15:0] apply_selecter_3_io_xbar_in_bits_tkeep; // @[BFS.scala 268:11]
  wire  apply_selecter_3_io_xbar_in_bits_tlast; // @[BFS.scala 268:11]
  wire  apply_selecter_3_io_ddr_out_ready; // @[BFS.scala 268:11]
  wire  apply_selecter_3_io_ddr_out_valid; // @[BFS.scala 268:11]
  wire [31:0] apply_selecter_3_io_ddr_out_bits_tdata; // @[BFS.scala 268:11]
  wire  vertex_update_buffer_0_full; // @[BFS.scala 271:11]
  wire [63:0] vertex_update_buffer_0_din; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_0_wr_en; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_0_empty; // @[BFS.scala 271:11]
  wire [63:0] vertex_update_buffer_0_dout; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_0_rd_en; // @[BFS.scala 271:11]
  wire [5:0] vertex_update_buffer_0_data_count; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_0_clk; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_0_srst; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_0_valid; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_1_full; // @[BFS.scala 271:11]
  wire [63:0] vertex_update_buffer_1_din; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_1_wr_en; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_1_empty; // @[BFS.scala 271:11]
  wire [63:0] vertex_update_buffer_1_dout; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_1_rd_en; // @[BFS.scala 271:11]
  wire [5:0] vertex_update_buffer_1_data_count; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_1_clk; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_1_srst; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_1_valid; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_2_full; // @[BFS.scala 271:11]
  wire [63:0] vertex_update_buffer_2_din; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_2_wr_en; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_2_empty; // @[BFS.scala 271:11]
  wire [63:0] vertex_update_buffer_2_dout; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_2_rd_en; // @[BFS.scala 271:11]
  wire [5:0] vertex_update_buffer_2_data_count; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_2_clk; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_2_srst; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_2_valid; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_3_full; // @[BFS.scala 271:11]
  wire [63:0] vertex_update_buffer_3_din; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_3_wr_en; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_3_empty; // @[BFS.scala 271:11]
  wire [63:0] vertex_update_buffer_3_dout; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_3_rd_en; // @[BFS.scala 271:11]
  wire [5:0] vertex_update_buffer_3_data_count; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_3_clk; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_3_srst; // @[BFS.scala 271:11]
  wire  vertex_update_buffer_3_valid; // @[BFS.scala 271:11]
  wire  update_engine_0_clock; // @[BFS.scala 274:16]
  wire  update_engine_0_reset; // @[BFS.scala 274:16]
  wire  update_engine_0_io_axi_ddr_aw_ready; // @[BFS.scala 274:16]
  wire  update_engine_0_io_axi_ddr_aw_valid; // @[BFS.scala 274:16]
  wire [63:0] update_engine_0_io_axi_ddr_aw_bits_awaddr; // @[BFS.scala 274:16]
  wire [5:0] update_engine_0_io_axi_ddr_aw_bits_awid; // @[BFS.scala 274:16]
  wire  update_engine_0_io_axi_ddr_w_ready; // @[BFS.scala 274:16]
  wire  update_engine_0_io_axi_ddr_w_valid; // @[BFS.scala 274:16]
  wire [127:0] update_engine_0_io_axi_ddr_w_bits_wdata; // @[BFS.scala 274:16]
  wire [15:0] update_engine_0_io_axi_ddr_w_bits_wstrb; // @[BFS.scala 274:16]
  wire  update_engine_0_io_xbar_in_ready; // @[BFS.scala 274:16]
  wire  update_engine_0_io_xbar_in_valid; // @[BFS.scala 274:16]
  wire [31:0] update_engine_0_io_xbar_in_bits_tdata; // @[BFS.scala 274:16]
  wire [63:0] update_engine_0_io_level_base_addr; // @[BFS.scala 274:16]
  wire [31:0] update_engine_0_io_level; // @[BFS.scala 274:16]
  wire  update_engine_0_io_end; // @[BFS.scala 274:16]
  wire  update_engine_0_io_flush; // @[BFS.scala 274:16]
  wire  update_engine_1_clock; // @[BFS.scala 274:16]
  wire  update_engine_1_reset; // @[BFS.scala 274:16]
  wire  update_engine_1_io_axi_ddr_aw_ready; // @[BFS.scala 274:16]
  wire  update_engine_1_io_axi_ddr_aw_valid; // @[BFS.scala 274:16]
  wire [63:0] update_engine_1_io_axi_ddr_aw_bits_awaddr; // @[BFS.scala 274:16]
  wire [5:0] update_engine_1_io_axi_ddr_aw_bits_awid; // @[BFS.scala 274:16]
  wire  update_engine_1_io_axi_ddr_w_ready; // @[BFS.scala 274:16]
  wire  update_engine_1_io_axi_ddr_w_valid; // @[BFS.scala 274:16]
  wire [127:0] update_engine_1_io_axi_ddr_w_bits_wdata; // @[BFS.scala 274:16]
  wire [15:0] update_engine_1_io_axi_ddr_w_bits_wstrb; // @[BFS.scala 274:16]
  wire  update_engine_1_io_xbar_in_ready; // @[BFS.scala 274:16]
  wire  update_engine_1_io_xbar_in_valid; // @[BFS.scala 274:16]
  wire [31:0] update_engine_1_io_xbar_in_bits_tdata; // @[BFS.scala 274:16]
  wire [63:0] update_engine_1_io_level_base_addr; // @[BFS.scala 274:16]
  wire [31:0] update_engine_1_io_level; // @[BFS.scala 274:16]
  wire  update_engine_1_io_end; // @[BFS.scala 274:16]
  wire  update_engine_1_io_flush; // @[BFS.scala 274:16]
  wire  update_engine_2_clock; // @[BFS.scala 274:16]
  wire  update_engine_2_reset; // @[BFS.scala 274:16]
  wire  update_engine_2_io_axi_ddr_aw_ready; // @[BFS.scala 274:16]
  wire  update_engine_2_io_axi_ddr_aw_valid; // @[BFS.scala 274:16]
  wire [63:0] update_engine_2_io_axi_ddr_aw_bits_awaddr; // @[BFS.scala 274:16]
  wire [5:0] update_engine_2_io_axi_ddr_aw_bits_awid; // @[BFS.scala 274:16]
  wire  update_engine_2_io_axi_ddr_w_ready; // @[BFS.scala 274:16]
  wire  update_engine_2_io_axi_ddr_w_valid; // @[BFS.scala 274:16]
  wire [127:0] update_engine_2_io_axi_ddr_w_bits_wdata; // @[BFS.scala 274:16]
  wire [15:0] update_engine_2_io_axi_ddr_w_bits_wstrb; // @[BFS.scala 274:16]
  wire  update_engine_2_io_xbar_in_ready; // @[BFS.scala 274:16]
  wire  update_engine_2_io_xbar_in_valid; // @[BFS.scala 274:16]
  wire [31:0] update_engine_2_io_xbar_in_bits_tdata; // @[BFS.scala 274:16]
  wire [63:0] update_engine_2_io_level_base_addr; // @[BFS.scala 274:16]
  wire [31:0] update_engine_2_io_level; // @[BFS.scala 274:16]
  wire  update_engine_2_io_end; // @[BFS.scala 274:16]
  wire  update_engine_2_io_flush; // @[BFS.scala 274:16]
  wire  update_engine_3_clock; // @[BFS.scala 274:16]
  wire  update_engine_3_reset; // @[BFS.scala 274:16]
  wire  update_engine_3_io_axi_ddr_aw_ready; // @[BFS.scala 274:16]
  wire  update_engine_3_io_axi_ddr_aw_valid; // @[BFS.scala 274:16]
  wire [63:0] update_engine_3_io_axi_ddr_aw_bits_awaddr; // @[BFS.scala 274:16]
  wire [5:0] update_engine_3_io_axi_ddr_aw_bits_awid; // @[BFS.scala 274:16]
  wire  update_engine_3_io_axi_ddr_w_ready; // @[BFS.scala 274:16]
  wire  update_engine_3_io_axi_ddr_w_valid; // @[BFS.scala 274:16]
  wire [127:0] update_engine_3_io_axi_ddr_w_bits_wdata; // @[BFS.scala 274:16]
  wire [15:0] update_engine_3_io_axi_ddr_w_bits_wstrb; // @[BFS.scala 274:16]
  wire  update_engine_3_io_xbar_in_ready; // @[BFS.scala 274:16]
  wire  update_engine_3_io_xbar_in_valid; // @[BFS.scala 274:16]
  wire [31:0] update_engine_3_io_xbar_in_bits_tdata; // @[BFS.scala 274:16]
  wire [63:0] update_engine_3_io_level_base_addr; // @[BFS.scala 274:16]
  wire [31:0] update_engine_3_io_level; // @[BFS.scala 274:16]
  wire  update_engine_3_io_end; // @[BFS.scala 274:16]
  wire  update_engine_3_io_flush; // @[BFS.scala 274:16]
    (*dont_touch = "true" *)reg [31:0] ready_counter; // @[BFS.scala 241:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 244:36]
  reg  end_reg_0; // @[BFS.scala 276:24]
  reg  end_reg_1; // @[BFS.scala 276:24]
  reg  end_reg_2; // @[BFS.scala 276:24]
  reg  end_reg_3; // @[BFS.scala 276:24]
  wire  _apply_selecter_0_io_xbar_in_valid_T_1 = apply_selecter_0_io_xbar_in_bits_tkeep != 16'h0; // @[BFS.scala 280:49]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_6 = ~broadcaster_m_axis_tdata[31] & broadcaster_m_axis_tdata[1:0] == 2'h0
    ; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_7 = broadcaster_m_axis_tkeep[0] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_6; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_14 = ~broadcaster_m_axis_tdata[63] & broadcaster_m_axis_tdata[33:32]
     == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_15 = broadcaster_m_axis_tkeep[1] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_14; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_22 = ~broadcaster_m_axis_tdata[95] & broadcaster_m_axis_tdata[65:64]
     == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_23 = broadcaster_m_axis_tkeep[2] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_22; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_30 = ~broadcaster_m_axis_tdata[127] & broadcaster_m_axis_tdata[97:96]
     == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_31 = broadcaster_m_axis_tkeep[3] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_30; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_38 = ~broadcaster_m_axis_tdata[159] & broadcaster_m_axis_tdata[129:128
    ] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_39 = broadcaster_m_axis_tkeep[4] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_38; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_46 = ~broadcaster_m_axis_tdata[191] & broadcaster_m_axis_tdata[161:160
    ] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_47 = broadcaster_m_axis_tkeep[5] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_46; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_54 = ~broadcaster_m_axis_tdata[223] & broadcaster_m_axis_tdata[193:192
    ] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_55 = broadcaster_m_axis_tkeep[6] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_54; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_62 = ~broadcaster_m_axis_tdata[255] & broadcaster_m_axis_tdata[225:224
    ] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_63 = broadcaster_m_axis_tkeep[7] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_62; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_70 = ~broadcaster_m_axis_tdata[287] & broadcaster_m_axis_tdata[257:256
    ] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_71 = broadcaster_m_axis_tkeep[8] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_70; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_78 = ~broadcaster_m_axis_tdata[319] & broadcaster_m_axis_tdata[289:288
    ] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_79 = broadcaster_m_axis_tkeep[9] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_78; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_86 = ~broadcaster_m_axis_tdata[351] & broadcaster_m_axis_tdata[321:320
    ] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_87 = broadcaster_m_axis_tkeep[10] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_86; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_94 = ~broadcaster_m_axis_tdata[383] & broadcaster_m_axis_tdata[353:352
    ] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_95 = broadcaster_m_axis_tkeep[11] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_94; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_102 = ~broadcaster_m_axis_tdata[415] & broadcaster_m_axis_tdata[385:
    384] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_103 = broadcaster_m_axis_tkeep[12] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_102; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_110 = ~broadcaster_m_axis_tdata[447] & broadcaster_m_axis_tdata[417:
    416] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_111 = broadcaster_m_axis_tkeep[13] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_110; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_118 = ~broadcaster_m_axis_tdata[479] & broadcaster_m_axis_tdata[449:
    448] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_119 = broadcaster_m_axis_tkeep[14] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_118; // @[BFS.scala 286:63]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_126 = ~broadcaster_m_axis_tdata[511] & broadcaster_m_axis_tdata[481:
    480] == 2'h0; // @[BFS.scala 248:21]
  wire  _apply_selecter_0_io_xbar_in_bits_tkeep_T_127 = broadcaster_m_axis_tkeep[15] &
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_126; // @[BFS.scala 286:63]
  wire [7:0] apply_selecter_0_io_xbar_in_bits_tkeep_lo = {_apply_selecter_0_io_xbar_in_bits_tkeep_T_63,
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_55,_apply_selecter_0_io_xbar_in_bits_tkeep_T_47,
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_39,_apply_selecter_0_io_xbar_in_bits_tkeep_T_31,
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_23,_apply_selecter_0_io_xbar_in_bits_tkeep_T_15,
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_7}; // @[BFS.scala 290:15]
  wire [7:0] apply_selecter_0_io_xbar_in_bits_tkeep_hi = {_apply_selecter_0_io_xbar_in_bits_tkeep_T_127,
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_119,_apply_selecter_0_io_xbar_in_bits_tkeep_T_111,
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_103,_apply_selecter_0_io_xbar_in_bits_tkeep_T_95,
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_87,_apply_selecter_0_io_xbar_in_bits_tkeep_T_79,
    _apply_selecter_0_io_xbar_in_bits_tkeep_T_71}; // @[BFS.scala 290:15]
  wire  _update_engine_0_io_flush_T = vertex_update_buffer_0_data_count == 6'h0; // @[util.scala 211:19]
  wire  _GEN_1 = update_engine_0_io_end | end_reg_0; // @[BFS.scala 307:36 BFS.scala 308:20 BFS.scala 276:24]
  wire  _apply_selecter_1_io_xbar_in_valid_T_1 = apply_selecter_1_io_xbar_in_bits_tkeep != 16'h0; // @[BFS.scala 280:49]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_6 = ~broadcaster_m_axis_tdata[543] & broadcaster_m_axis_tdata[513:512]
     == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_7 = broadcaster_m_axis_tkeep[64] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_6; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_14 = ~broadcaster_m_axis_tdata[575] & broadcaster_m_axis_tdata[545:544
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_15 = broadcaster_m_axis_tkeep[65] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_14; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_22 = ~broadcaster_m_axis_tdata[607] & broadcaster_m_axis_tdata[577:576
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_23 = broadcaster_m_axis_tkeep[66] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_22; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_30 = ~broadcaster_m_axis_tdata[639] & broadcaster_m_axis_tdata[609:608
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_31 = broadcaster_m_axis_tkeep[67] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_30; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_38 = ~broadcaster_m_axis_tdata[671] & broadcaster_m_axis_tdata[641:640
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_39 = broadcaster_m_axis_tkeep[68] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_38; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_46 = ~broadcaster_m_axis_tdata[703] & broadcaster_m_axis_tdata[673:672
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_47 = broadcaster_m_axis_tkeep[69] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_46; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_54 = ~broadcaster_m_axis_tdata[735] & broadcaster_m_axis_tdata[705:704
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_55 = broadcaster_m_axis_tkeep[70] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_54; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_62 = ~broadcaster_m_axis_tdata[767] & broadcaster_m_axis_tdata[737:736
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_63 = broadcaster_m_axis_tkeep[71] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_62; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_70 = ~broadcaster_m_axis_tdata[799] & broadcaster_m_axis_tdata[769:768
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_71 = broadcaster_m_axis_tkeep[72] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_70; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_78 = ~broadcaster_m_axis_tdata[831] & broadcaster_m_axis_tdata[801:800
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_79 = broadcaster_m_axis_tkeep[73] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_78; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_86 = ~broadcaster_m_axis_tdata[863] & broadcaster_m_axis_tdata[833:832
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_87 = broadcaster_m_axis_tkeep[74] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_86; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_94 = ~broadcaster_m_axis_tdata[895] & broadcaster_m_axis_tdata[865:864
    ] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_95 = broadcaster_m_axis_tkeep[75] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_94; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_102 = ~broadcaster_m_axis_tdata[927] & broadcaster_m_axis_tdata[897:
    896] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_103 = broadcaster_m_axis_tkeep[76] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_102; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_110 = ~broadcaster_m_axis_tdata[959] & broadcaster_m_axis_tdata[929:
    928] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_111 = broadcaster_m_axis_tkeep[77] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_110; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_118 = ~broadcaster_m_axis_tdata[991] & broadcaster_m_axis_tdata[961:
    960] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_119 = broadcaster_m_axis_tkeep[78] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_118; // @[BFS.scala 286:63]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_126 = ~broadcaster_m_axis_tdata[1023] & broadcaster_m_axis_tdata[993:
    992] == 2'h1; // @[BFS.scala 248:21]
  wire  _apply_selecter_1_io_xbar_in_bits_tkeep_T_127 = broadcaster_m_axis_tkeep[79] &
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_126; // @[BFS.scala 286:63]
  wire [7:0] apply_selecter_1_io_xbar_in_bits_tkeep_lo = {_apply_selecter_1_io_xbar_in_bits_tkeep_T_63,
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_55,_apply_selecter_1_io_xbar_in_bits_tkeep_T_47,
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_39,_apply_selecter_1_io_xbar_in_bits_tkeep_T_31,
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_23,_apply_selecter_1_io_xbar_in_bits_tkeep_T_15,
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_7}; // @[BFS.scala 290:15]
  wire [7:0] apply_selecter_1_io_xbar_in_bits_tkeep_hi = {_apply_selecter_1_io_xbar_in_bits_tkeep_T_127,
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_119,_apply_selecter_1_io_xbar_in_bits_tkeep_T_111,
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_103,_apply_selecter_1_io_xbar_in_bits_tkeep_T_95,
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_87,_apply_selecter_1_io_xbar_in_bits_tkeep_T_79,
    _apply_selecter_1_io_xbar_in_bits_tkeep_T_71}; // @[BFS.scala 290:15]
  wire  _update_engine_1_io_flush_T = vertex_update_buffer_1_data_count == 6'h0; // @[util.scala 211:19]
  wire  _GEN_2 = update_engine_1_io_end | end_reg_1; // @[BFS.scala 307:36 BFS.scala 308:20 BFS.scala 276:24]
  wire  _apply_selecter_2_io_xbar_in_valid_T_1 = apply_selecter_2_io_xbar_in_bits_tkeep != 16'h0; // @[BFS.scala 280:49]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_6 = ~broadcaster_m_axis_tdata[1055] & broadcaster_m_axis_tdata[1025:
    1024] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_7 = broadcaster_m_axis_tkeep[128] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_6; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_14 = ~broadcaster_m_axis_tdata[1087] & broadcaster_m_axis_tdata[1057:
    1056] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_15 = broadcaster_m_axis_tkeep[129] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_14; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_22 = ~broadcaster_m_axis_tdata[1119] & broadcaster_m_axis_tdata[1089:
    1088] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_23 = broadcaster_m_axis_tkeep[130] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_22; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_30 = ~broadcaster_m_axis_tdata[1151] & broadcaster_m_axis_tdata[1121:
    1120] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_31 = broadcaster_m_axis_tkeep[131] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_30; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_38 = ~broadcaster_m_axis_tdata[1183] & broadcaster_m_axis_tdata[1153:
    1152] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_39 = broadcaster_m_axis_tkeep[132] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_38; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_46 = ~broadcaster_m_axis_tdata[1215] & broadcaster_m_axis_tdata[1185:
    1184] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_47 = broadcaster_m_axis_tkeep[133] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_46; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_54 = ~broadcaster_m_axis_tdata[1247] & broadcaster_m_axis_tdata[1217:
    1216] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_55 = broadcaster_m_axis_tkeep[134] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_54; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_62 = ~broadcaster_m_axis_tdata[1279] & broadcaster_m_axis_tdata[1249:
    1248] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_63 = broadcaster_m_axis_tkeep[135] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_62; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_70 = ~broadcaster_m_axis_tdata[1311] & broadcaster_m_axis_tdata[1281:
    1280] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_71 = broadcaster_m_axis_tkeep[136] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_70; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_78 = ~broadcaster_m_axis_tdata[1343] & broadcaster_m_axis_tdata[1313:
    1312] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_79 = broadcaster_m_axis_tkeep[137] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_78; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_86 = ~broadcaster_m_axis_tdata[1375] & broadcaster_m_axis_tdata[1345:
    1344] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_87 = broadcaster_m_axis_tkeep[138] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_86; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_94 = ~broadcaster_m_axis_tdata[1407] & broadcaster_m_axis_tdata[1377:
    1376] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_95 = broadcaster_m_axis_tkeep[139] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_94; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_102 = ~broadcaster_m_axis_tdata[1439] & broadcaster_m_axis_tdata[1409:
    1408] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_103 = broadcaster_m_axis_tkeep[140] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_102; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_110 = ~broadcaster_m_axis_tdata[1471] & broadcaster_m_axis_tdata[1441:
    1440] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_111 = broadcaster_m_axis_tkeep[141] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_110; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_118 = ~broadcaster_m_axis_tdata[1503] & broadcaster_m_axis_tdata[1473:
    1472] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_119 = broadcaster_m_axis_tkeep[142] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_118; // @[BFS.scala 286:63]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_126 = ~broadcaster_m_axis_tdata[1535] & broadcaster_m_axis_tdata[1505:
    1504] == 2'h2; // @[BFS.scala 248:21]
  wire  _apply_selecter_2_io_xbar_in_bits_tkeep_T_127 = broadcaster_m_axis_tkeep[143] &
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_126; // @[BFS.scala 286:63]
  wire [7:0] apply_selecter_2_io_xbar_in_bits_tkeep_lo = {_apply_selecter_2_io_xbar_in_bits_tkeep_T_63,
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_55,_apply_selecter_2_io_xbar_in_bits_tkeep_T_47,
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_39,_apply_selecter_2_io_xbar_in_bits_tkeep_T_31,
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_23,_apply_selecter_2_io_xbar_in_bits_tkeep_T_15,
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_7}; // @[BFS.scala 290:15]
  wire [7:0] apply_selecter_2_io_xbar_in_bits_tkeep_hi = {_apply_selecter_2_io_xbar_in_bits_tkeep_T_127,
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_119,_apply_selecter_2_io_xbar_in_bits_tkeep_T_111,
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_103,_apply_selecter_2_io_xbar_in_bits_tkeep_T_95,
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_87,_apply_selecter_2_io_xbar_in_bits_tkeep_T_79,
    _apply_selecter_2_io_xbar_in_bits_tkeep_T_71}; // @[BFS.scala 290:15]
  wire  _update_engine_2_io_flush_T = vertex_update_buffer_2_data_count == 6'h0; // @[util.scala 211:19]
  wire  _GEN_3 = update_engine_2_io_end | end_reg_2; // @[BFS.scala 307:36 BFS.scala 308:20 BFS.scala 276:24]
  wire  _apply_selecter_3_io_xbar_in_valid_T_1 = apply_selecter_3_io_xbar_in_bits_tkeep != 16'h0; // @[BFS.scala 280:49]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_6 = ~broadcaster_m_axis_tdata[1567] & broadcaster_m_axis_tdata[1537:
    1536] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_7 = broadcaster_m_axis_tkeep[192] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_6; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_14 = ~broadcaster_m_axis_tdata[1599] & broadcaster_m_axis_tdata[1569:
    1568] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_15 = broadcaster_m_axis_tkeep[193] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_14; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_22 = ~broadcaster_m_axis_tdata[1631] & broadcaster_m_axis_tdata[1601:
    1600] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_23 = broadcaster_m_axis_tkeep[194] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_22; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_30 = ~broadcaster_m_axis_tdata[1663] & broadcaster_m_axis_tdata[1633:
    1632] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_31 = broadcaster_m_axis_tkeep[195] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_30; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_38 = ~broadcaster_m_axis_tdata[1695] & broadcaster_m_axis_tdata[1665:
    1664] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_39 = broadcaster_m_axis_tkeep[196] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_38; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_46 = ~broadcaster_m_axis_tdata[1727] & broadcaster_m_axis_tdata[1697:
    1696] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_47 = broadcaster_m_axis_tkeep[197] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_46; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_54 = ~broadcaster_m_axis_tdata[1759] & broadcaster_m_axis_tdata[1729:
    1728] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_55 = broadcaster_m_axis_tkeep[198] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_54; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_62 = ~broadcaster_m_axis_tdata[1791] & broadcaster_m_axis_tdata[1761:
    1760] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_63 = broadcaster_m_axis_tkeep[199] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_62; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_70 = ~broadcaster_m_axis_tdata[1823] & broadcaster_m_axis_tdata[1793:
    1792] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_71 = broadcaster_m_axis_tkeep[200] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_70; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_78 = ~broadcaster_m_axis_tdata[1855] & broadcaster_m_axis_tdata[1825:
    1824] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_79 = broadcaster_m_axis_tkeep[201] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_78; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_86 = ~broadcaster_m_axis_tdata[1887] & broadcaster_m_axis_tdata[1857:
    1856] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_87 = broadcaster_m_axis_tkeep[202] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_86; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_94 = ~broadcaster_m_axis_tdata[1919] & broadcaster_m_axis_tdata[1889:
    1888] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_95 = broadcaster_m_axis_tkeep[203] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_94; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_102 = ~broadcaster_m_axis_tdata[1951] & broadcaster_m_axis_tdata[1921:
    1920] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_103 = broadcaster_m_axis_tkeep[204] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_102; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_110 = ~broadcaster_m_axis_tdata[1983] & broadcaster_m_axis_tdata[1953:
    1952] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_111 = broadcaster_m_axis_tkeep[205] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_110; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_118 = ~broadcaster_m_axis_tdata[2015] & broadcaster_m_axis_tdata[1985:
    1984] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_119 = broadcaster_m_axis_tkeep[206] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_118; // @[BFS.scala 286:63]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_126 = ~broadcaster_m_axis_tdata[2047] & broadcaster_m_axis_tdata[2017:
    2016] == 2'h3; // @[BFS.scala 248:21]
  wire  _apply_selecter_3_io_xbar_in_bits_tkeep_T_127 = broadcaster_m_axis_tkeep[207] &
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_126; // @[BFS.scala 286:63]
  wire [7:0] apply_selecter_3_io_xbar_in_bits_tkeep_lo = {_apply_selecter_3_io_xbar_in_bits_tkeep_T_63,
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_55,_apply_selecter_3_io_xbar_in_bits_tkeep_T_47,
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_39,_apply_selecter_3_io_xbar_in_bits_tkeep_T_31,
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_23,_apply_selecter_3_io_xbar_in_bits_tkeep_T_15,
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_7}; // @[BFS.scala 290:15]
  wire [7:0] apply_selecter_3_io_xbar_in_bits_tkeep_hi = {_apply_selecter_3_io_xbar_in_bits_tkeep_T_127,
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_119,_apply_selecter_3_io_xbar_in_bits_tkeep_T_111,
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_103,_apply_selecter_3_io_xbar_in_bits_tkeep_T_95,
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_87,_apply_selecter_3_io_xbar_in_bits_tkeep_T_79,
    _apply_selecter_3_io_xbar_in_bits_tkeep_T_71}; // @[BFS.scala 290:15]
  wire  _update_engine_3_io_flush_T = vertex_update_buffer_3_data_count == 6'h0; // @[util.scala 211:19]
  wire  _GEN_4 = update_engine_3_io_end | end_reg_3; // @[BFS.scala 307:36 BFS.scala 308:20 BFS.scala 276:24]
  wire  _broadcaster_io_m_axis_tready_WIRE_1 = apply_selecter_1_io_xbar_in_ready; // @[BFS.scala 312:42 BFS.scala 312:42]
  wire  _broadcaster_io_m_axis_tready_WIRE_0 = apply_selecter_0_io_xbar_in_ready; // @[BFS.scala 312:42 BFS.scala 312:42]
  wire [1:0] broadcaster_io_m_axis_tready_lo = {_broadcaster_io_m_axis_tready_WIRE_1,
    _broadcaster_io_m_axis_tready_WIRE_0}; // @[BFS.scala 312:92]
  wire  _broadcaster_io_m_axis_tready_WIRE_3 = apply_selecter_3_io_xbar_in_ready; // @[BFS.scala 312:42 BFS.scala 312:42]
  wire  _broadcaster_io_m_axis_tready_WIRE_2 = apply_selecter_2_io_xbar_in_ready; // @[BFS.scala 312:42 BFS.scala 312:42]
  wire [1:0] broadcaster_io_m_axis_tready_hi = {_broadcaster_io_m_axis_tready_WIRE_3,
    _broadcaster_io_m_axis_tready_WIRE_2}; // @[BFS.scala 312:92]
  v2A_reg_slice apply_in ( // @[BFS.scala 251:24]
    .aclk(apply_in_aclk),
    .aresetn(apply_in_aresetn),
    .s_axis_tdata(apply_in_s_axis_tdata),
    .s_axis_tkeep(apply_in_s_axis_tkeep),
    .s_axis_tvalid(apply_in_s_axis_tvalid),
    .s_axis_tready(apply_in_s_axis_tready),
    .s_axis_tlast(apply_in_s_axis_tlast),
    .m_axis_tdata(apply_in_m_axis_tdata),
    .m_axis_tkeep(apply_in_m_axis_tkeep),
    .m_axis_tvalid(apply_in_m_axis_tvalid),
    .m_axis_tready(apply_in_m_axis_tready),
    .m_axis_tlast(apply_in_m_axis_tlast)
  );
  level_cache_broadcaster broadcaster ( // @[BFS.scala 258:27]
    .aclk(broadcaster_aclk),
    .aresetn(broadcaster_aresetn),
    .s_axis_tdata(broadcaster_s_axis_tdata),
    .s_axis_tkeep(broadcaster_s_axis_tkeep),
    .s_axis_tvalid(broadcaster_s_axis_tvalid),
    .s_axis_tready(broadcaster_s_axis_tready),
    .s_axis_tlast(broadcaster_s_axis_tlast),
    .s_axis_tid(broadcaster_s_axis_tid),
    .m_axis_tdata(broadcaster_m_axis_tdata),
    .m_axis_tkeep(broadcaster_m_axis_tkeep),
    .m_axis_tvalid(broadcaster_m_axis_tvalid),
    .m_axis_tready(broadcaster_m_axis_tready),
    .m_axis_tlast(broadcaster_m_axis_tlast),
    .m_axis_tid(broadcaster_m_axis_tid)
  );
  axis_arbitrator apply_selecter_0 ( // @[BFS.scala 268:11]
    .clock(apply_selecter_0_clock),
    .reset(apply_selecter_0_reset),
    .io_xbar_in_ready(apply_selecter_0_io_xbar_in_ready),
    .io_xbar_in_valid(apply_selecter_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(apply_selecter_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(apply_selecter_0_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(apply_selecter_0_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(apply_selecter_0_io_ddr_out_ready),
    .io_ddr_out_valid(apply_selecter_0_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(apply_selecter_0_io_ddr_out_bits_tdata)
  );
  axis_arbitrator apply_selecter_1 ( // @[BFS.scala 268:11]
    .clock(apply_selecter_1_clock),
    .reset(apply_selecter_1_reset),
    .io_xbar_in_ready(apply_selecter_1_io_xbar_in_ready),
    .io_xbar_in_valid(apply_selecter_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(apply_selecter_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(apply_selecter_1_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(apply_selecter_1_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(apply_selecter_1_io_ddr_out_ready),
    .io_ddr_out_valid(apply_selecter_1_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(apply_selecter_1_io_ddr_out_bits_tdata)
  );
  axis_arbitrator apply_selecter_2 ( // @[BFS.scala 268:11]
    .clock(apply_selecter_2_clock),
    .reset(apply_selecter_2_reset),
    .io_xbar_in_ready(apply_selecter_2_io_xbar_in_ready),
    .io_xbar_in_valid(apply_selecter_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(apply_selecter_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(apply_selecter_2_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(apply_selecter_2_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(apply_selecter_2_io_ddr_out_ready),
    .io_ddr_out_valid(apply_selecter_2_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(apply_selecter_2_io_ddr_out_bits_tdata)
  );
  axis_arbitrator apply_selecter_3 ( // @[BFS.scala 268:11]
    .clock(apply_selecter_3_clock),
    .reset(apply_selecter_3_reset),
    .io_xbar_in_ready(apply_selecter_3_io_xbar_in_ready),
    .io_xbar_in_valid(apply_selecter_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(apply_selecter_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(apply_selecter_3_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(apply_selecter_3_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(apply_selecter_3_io_ddr_out_ready),
    .io_ddr_out_valid(apply_selecter_3_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(apply_selecter_3_io_ddr_out_bits_tdata)
  );
  update_fifo vertex_update_buffer_0 ( // @[BFS.scala 271:11]
    .full(vertex_update_buffer_0_full),
    .din(vertex_update_buffer_0_din),
    .wr_en(vertex_update_buffer_0_wr_en),
    .empty(vertex_update_buffer_0_empty),
    .dout(vertex_update_buffer_0_dout),
    .rd_en(vertex_update_buffer_0_rd_en),
    .data_count(vertex_update_buffer_0_data_count),
    .clk(vertex_update_buffer_0_clk),
    .srst(vertex_update_buffer_0_srst),
    .valid(vertex_update_buffer_0_valid)
  );
  update_fifo vertex_update_buffer_1 ( // @[BFS.scala 271:11]
    .full(vertex_update_buffer_1_full),
    .din(vertex_update_buffer_1_din),
    .wr_en(vertex_update_buffer_1_wr_en),
    .empty(vertex_update_buffer_1_empty),
    .dout(vertex_update_buffer_1_dout),
    .rd_en(vertex_update_buffer_1_rd_en),
    .data_count(vertex_update_buffer_1_data_count),
    .clk(vertex_update_buffer_1_clk),
    .srst(vertex_update_buffer_1_srst),
    .valid(vertex_update_buffer_1_valid)
  );
  update_fifo vertex_update_buffer_2 ( // @[BFS.scala 271:11]
    .full(vertex_update_buffer_2_full),
    .din(vertex_update_buffer_2_din),
    .wr_en(vertex_update_buffer_2_wr_en),
    .empty(vertex_update_buffer_2_empty),
    .dout(vertex_update_buffer_2_dout),
    .rd_en(vertex_update_buffer_2_rd_en),
    .data_count(vertex_update_buffer_2_data_count),
    .clk(vertex_update_buffer_2_clk),
    .srst(vertex_update_buffer_2_srst),
    .valid(vertex_update_buffer_2_valid)
  );
  update_fifo vertex_update_buffer_3 ( // @[BFS.scala 271:11]
    .full(vertex_update_buffer_3_full),
    .din(vertex_update_buffer_3_din),
    .wr_en(vertex_update_buffer_3_wr_en),
    .empty(vertex_update_buffer_3_empty),
    .dout(vertex_update_buffer_3_dout),
    .rd_en(vertex_update_buffer_3_rd_en),
    .data_count(vertex_update_buffer_3_data_count),
    .clk(vertex_update_buffer_3_clk),
    .srst(vertex_update_buffer_3_srst),
    .valid(vertex_update_buffer_3_valid)
  );
  WB_engine update_engine_0 ( // @[BFS.scala 274:16]
    .clock(update_engine_0_clock),
    .reset(update_engine_0_reset),
    .io_axi_ddr_aw_ready(update_engine_0_io_axi_ddr_aw_ready),
    .io_axi_ddr_aw_valid(update_engine_0_io_axi_ddr_aw_valid),
    .io_axi_ddr_aw_bits_awaddr(update_engine_0_io_axi_ddr_aw_bits_awaddr),
    .io_axi_ddr_aw_bits_awid(update_engine_0_io_axi_ddr_aw_bits_awid),
    .io_axi_ddr_w_ready(update_engine_0_io_axi_ddr_w_ready),
    .io_axi_ddr_w_valid(update_engine_0_io_axi_ddr_w_valid),
    .io_axi_ddr_w_bits_wdata(update_engine_0_io_axi_ddr_w_bits_wdata),
    .io_axi_ddr_w_bits_wstrb(update_engine_0_io_axi_ddr_w_bits_wstrb),
    .io_xbar_in_ready(update_engine_0_io_xbar_in_ready),
    .io_xbar_in_valid(update_engine_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(update_engine_0_io_xbar_in_bits_tdata),
    .io_level_base_addr(update_engine_0_io_level_base_addr),
    .io_level(update_engine_0_io_level),
    .io_end(update_engine_0_io_end),
    .io_flush(update_engine_0_io_flush)
  );
  WB_engine_1 update_engine_1 ( // @[BFS.scala 274:16]
    .clock(update_engine_1_clock),
    .reset(update_engine_1_reset),
    .io_axi_ddr_aw_ready(update_engine_1_io_axi_ddr_aw_ready),
    .io_axi_ddr_aw_valid(update_engine_1_io_axi_ddr_aw_valid),
    .io_axi_ddr_aw_bits_awaddr(update_engine_1_io_axi_ddr_aw_bits_awaddr),
    .io_axi_ddr_aw_bits_awid(update_engine_1_io_axi_ddr_aw_bits_awid),
    .io_axi_ddr_w_ready(update_engine_1_io_axi_ddr_w_ready),
    .io_axi_ddr_w_valid(update_engine_1_io_axi_ddr_w_valid),
    .io_axi_ddr_w_bits_wdata(update_engine_1_io_axi_ddr_w_bits_wdata),
    .io_axi_ddr_w_bits_wstrb(update_engine_1_io_axi_ddr_w_bits_wstrb),
    .io_xbar_in_ready(update_engine_1_io_xbar_in_ready),
    .io_xbar_in_valid(update_engine_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(update_engine_1_io_xbar_in_bits_tdata),
    .io_level_base_addr(update_engine_1_io_level_base_addr),
    .io_level(update_engine_1_io_level),
    .io_end(update_engine_1_io_end),
    .io_flush(update_engine_1_io_flush)
  );
  WB_engine_2 update_engine_2 ( // @[BFS.scala 274:16]
    .clock(update_engine_2_clock),
    .reset(update_engine_2_reset),
    .io_axi_ddr_aw_ready(update_engine_2_io_axi_ddr_aw_ready),
    .io_axi_ddr_aw_valid(update_engine_2_io_axi_ddr_aw_valid),
    .io_axi_ddr_aw_bits_awaddr(update_engine_2_io_axi_ddr_aw_bits_awaddr),
    .io_axi_ddr_aw_bits_awid(update_engine_2_io_axi_ddr_aw_bits_awid),
    .io_axi_ddr_w_ready(update_engine_2_io_axi_ddr_w_ready),
    .io_axi_ddr_w_valid(update_engine_2_io_axi_ddr_w_valid),
    .io_axi_ddr_w_bits_wdata(update_engine_2_io_axi_ddr_w_bits_wdata),
    .io_axi_ddr_w_bits_wstrb(update_engine_2_io_axi_ddr_w_bits_wstrb),
    .io_xbar_in_ready(update_engine_2_io_xbar_in_ready),
    .io_xbar_in_valid(update_engine_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(update_engine_2_io_xbar_in_bits_tdata),
    .io_level_base_addr(update_engine_2_io_level_base_addr),
    .io_level(update_engine_2_io_level),
    .io_end(update_engine_2_io_end),
    .io_flush(update_engine_2_io_flush)
  );
  WB_engine_3 update_engine_3 ( // @[BFS.scala 274:16]
    .clock(update_engine_3_clock),
    .reset(update_engine_3_reset),
    .io_axi_ddr_aw_ready(update_engine_3_io_axi_ddr_aw_ready),
    .io_axi_ddr_aw_valid(update_engine_3_io_axi_ddr_aw_valid),
    .io_axi_ddr_aw_bits_awaddr(update_engine_3_io_axi_ddr_aw_bits_awaddr),
    .io_axi_ddr_aw_bits_awid(update_engine_3_io_axi_ddr_aw_bits_awid),
    .io_axi_ddr_w_ready(update_engine_3_io_axi_ddr_w_ready),
    .io_axi_ddr_w_valid(update_engine_3_io_axi_ddr_w_valid),
    .io_axi_ddr_w_bits_wdata(update_engine_3_io_axi_ddr_w_bits_wdata),
    .io_axi_ddr_w_bits_wstrb(update_engine_3_io_axi_ddr_w_bits_wstrb),
    .io_xbar_in_ready(update_engine_3_io_xbar_in_ready),
    .io_xbar_in_valid(update_engine_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(update_engine_3_io_xbar_in_bits_tdata),
    .io_level_base_addr(update_engine_3_io_level_base_addr),
    .io_level(update_engine_3_io_level),
    .io_end(update_engine_3_io_end),
    .io_flush(update_engine_3_io_flush)
  );
  assign io_axi_0_ddr_aw_valid = update_engine_0_io_axi_ddr_aw_valid; // @[BFS.scala 305:17]
  assign io_axi_0_ddr_aw_bits_awaddr = update_engine_0_io_axi_ddr_aw_bits_awaddr; // @[BFS.scala 305:17]
  assign io_axi_0_ddr_aw_bits_awid = update_engine_0_io_axi_ddr_aw_bits_awid; // @[BFS.scala 305:17]
  assign io_axi_0_ddr_w_valid = update_engine_0_io_axi_ddr_w_valid; // @[BFS.scala 305:17]
  assign io_axi_0_ddr_w_bits_wdata = update_engine_0_io_axi_ddr_w_bits_wdata; // @[BFS.scala 305:17]
  assign io_axi_0_ddr_w_bits_wstrb = update_engine_0_io_axi_ddr_w_bits_wstrb; // @[BFS.scala 305:17]
  assign io_axi_1_ddr_aw_valid = update_engine_1_io_axi_ddr_aw_valid; // @[BFS.scala 305:17]
  assign io_axi_1_ddr_aw_bits_awaddr = update_engine_1_io_axi_ddr_aw_bits_awaddr; // @[BFS.scala 305:17]
  assign io_axi_1_ddr_aw_bits_awid = update_engine_1_io_axi_ddr_aw_bits_awid; // @[BFS.scala 305:17]
  assign io_axi_1_ddr_w_valid = update_engine_1_io_axi_ddr_w_valid; // @[BFS.scala 305:17]
  assign io_axi_1_ddr_w_bits_wdata = update_engine_1_io_axi_ddr_w_bits_wdata; // @[BFS.scala 305:17]
  assign io_axi_1_ddr_w_bits_wstrb = update_engine_1_io_axi_ddr_w_bits_wstrb; // @[BFS.scala 305:17]
  assign io_axi_2_ddr_aw_valid = update_engine_2_io_axi_ddr_aw_valid; // @[BFS.scala 305:17]
  assign io_axi_2_ddr_aw_bits_awaddr = update_engine_2_io_axi_ddr_aw_bits_awaddr; // @[BFS.scala 305:17]
  assign io_axi_2_ddr_aw_bits_awid = update_engine_2_io_axi_ddr_aw_bits_awid; // @[BFS.scala 305:17]
  assign io_axi_2_ddr_w_valid = update_engine_2_io_axi_ddr_w_valid; // @[BFS.scala 305:17]
  assign io_axi_2_ddr_w_bits_wdata = update_engine_2_io_axi_ddr_w_bits_wdata; // @[BFS.scala 305:17]
  assign io_axi_2_ddr_w_bits_wstrb = update_engine_2_io_axi_ddr_w_bits_wstrb; // @[BFS.scala 305:17]
  assign io_axi_3_ddr_aw_valid = update_engine_3_io_axi_ddr_aw_valid; // @[BFS.scala 305:17]
  assign io_axi_3_ddr_aw_bits_awaddr = update_engine_3_io_axi_ddr_aw_bits_awaddr; // @[BFS.scala 305:17]
  assign io_axi_3_ddr_aw_bits_awid = update_engine_3_io_axi_ddr_aw_bits_awid; // @[BFS.scala 305:17]
  assign io_axi_3_ddr_w_valid = update_engine_3_io_axi_ddr_w_valid; // @[BFS.scala 305:17]
  assign io_axi_3_ddr_w_bits_wdata = update_engine_3_io_axi_ddr_w_bits_wdata; // @[BFS.scala 305:17]
  assign io_axi_3_ddr_w_bits_wstrb = update_engine_3_io_axi_ddr_w_bits_wstrb; // @[BFS.scala 305:17]
  assign io_gather_in_ready = apply_in_s_axis_tready; // @[BFS.scala 256:22]
  assign io_end = end_reg_0 & end_reg_1 & end_reg_2 & end_reg_3; // @[BFS.scala 314:29]
  assign apply_in_aclk = clock; // @[BFS.scala 252:35]
  assign apply_in_aresetn = ~reset; // @[BFS.scala 253:26]
  assign apply_in_s_axis_tdata = io_gather_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign apply_in_s_axis_tkeep = io_gather_in_bits_tkeep; // @[nf_arm_doce_top.scala 121:11]
  assign apply_in_s_axis_tvalid = io_gather_in_valid; // @[BFS.scala 255:29]
  assign apply_in_s_axis_tlast = io_gather_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign apply_in_m_axis_tready = broadcaster_s_axis_tready; // @[BFS.scala 265:29]
  assign broadcaster_aclk = clock; // @[BFS.scala 260:38]
  assign broadcaster_aresetn = ~reset; // @[BFS.scala 259:29]
  assign broadcaster_s_axis_tdata = apply_in_m_axis_tdata; // @[BFS.scala 263:31]
  assign broadcaster_s_axis_tkeep = apply_in_m_axis_tkeep; // @[BFS.scala 262:31]
  assign broadcaster_s_axis_tvalid = apply_in_m_axis_tvalid; // @[BFS.scala 261:32]
  assign broadcaster_s_axis_tlast = apply_in_m_axis_tlast; // @[BFS.scala 264:31]
  assign broadcaster_s_axis_tid = 1'h0;
  assign broadcaster_m_axis_tready = {broadcaster_io_m_axis_tready_hi,broadcaster_io_m_axis_tready_lo}; // @[BFS.scala 312:92]
  assign apply_selecter_0_clock = clock;
  assign apply_selecter_0_reset = reset;
  assign apply_selecter_0_io_xbar_in_valid = broadcaster_m_axis_tvalid[0] & _apply_selecter_0_io_xbar_in_valid_T_1; // @[BFS.scala 279:77]
  assign apply_selecter_0_io_xbar_in_bits_tdata = broadcaster_m_axis_tdata[511:0]; // @[BFS.scala 283:36]
  assign apply_selecter_0_io_xbar_in_bits_tkeep = {apply_selecter_0_io_xbar_in_bits_tkeep_hi,
    apply_selecter_0_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 290:15]
  assign apply_selecter_0_io_xbar_in_bits_tlast = broadcaster_m_axis_tlast[0]; // @[BFS.scala 281:77]
  assign apply_selecter_0_io_ddr_out_ready = ~vertex_update_buffer_0_full; // @[util.scala 219:13]
  assign apply_selecter_1_clock = clock;
  assign apply_selecter_1_reset = reset;
  assign apply_selecter_1_io_xbar_in_valid = broadcaster_m_axis_tvalid[1] & _apply_selecter_1_io_xbar_in_valid_T_1; // @[BFS.scala 279:77]
  assign apply_selecter_1_io_xbar_in_bits_tdata = broadcaster_m_axis_tdata[1023:512]; // @[BFS.scala 283:36]
  assign apply_selecter_1_io_xbar_in_bits_tkeep = {apply_selecter_1_io_xbar_in_bits_tkeep_hi,
    apply_selecter_1_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 290:15]
  assign apply_selecter_1_io_xbar_in_bits_tlast = broadcaster_m_axis_tlast[1]; // @[BFS.scala 281:77]
  assign apply_selecter_1_io_ddr_out_ready = ~vertex_update_buffer_1_full; // @[util.scala 219:13]
  assign apply_selecter_2_clock = clock;
  assign apply_selecter_2_reset = reset;
  assign apply_selecter_2_io_xbar_in_valid = broadcaster_m_axis_tvalid[2] & _apply_selecter_2_io_xbar_in_valid_T_1; // @[BFS.scala 279:77]
  assign apply_selecter_2_io_xbar_in_bits_tdata = broadcaster_m_axis_tdata[1535:1024]; // @[BFS.scala 283:36]
  assign apply_selecter_2_io_xbar_in_bits_tkeep = {apply_selecter_2_io_xbar_in_bits_tkeep_hi,
    apply_selecter_2_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 290:15]
  assign apply_selecter_2_io_xbar_in_bits_tlast = broadcaster_m_axis_tlast[2]; // @[BFS.scala 281:77]
  assign apply_selecter_2_io_ddr_out_ready = ~vertex_update_buffer_2_full; // @[util.scala 219:13]
  assign apply_selecter_3_clock = clock;
  assign apply_selecter_3_reset = reset;
  assign apply_selecter_3_io_xbar_in_valid = broadcaster_m_axis_tvalid[3] & _apply_selecter_3_io_xbar_in_valid_T_1; // @[BFS.scala 279:77]
  assign apply_selecter_3_io_xbar_in_bits_tdata = broadcaster_m_axis_tdata[2047:1536]; // @[BFS.scala 283:36]
  assign apply_selecter_3_io_xbar_in_bits_tkeep = {apply_selecter_3_io_xbar_in_bits_tkeep_hi,
    apply_selecter_3_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 290:15]
  assign apply_selecter_3_io_xbar_in_bits_tlast = broadcaster_m_axis_tlast[3]; // @[BFS.scala 281:77]
  assign apply_selecter_3_io_ddr_out_ready = ~vertex_update_buffer_3_full; // @[util.scala 219:13]
  assign vertex_update_buffer_0_din = {apply_selecter_0_io_ddr_out_bits_tdata,io_level}; // @[Cat.scala 30:58]
  assign vertex_update_buffer_0_wr_en = apply_selecter_0_io_ddr_out_valid; // @[BFS.scala 294:40]
  assign vertex_update_buffer_0_rd_en = update_engine_0_io_xbar_in_ready; // @[BFS.scala 306:40]
  assign vertex_update_buffer_0_clk = clock; // @[BFS.scala 292:53]
  assign vertex_update_buffer_0_srst = reset; // @[BFS.scala 293:54]
  assign vertex_update_buffer_1_din = {apply_selecter_1_io_ddr_out_bits_tdata,io_level}; // @[Cat.scala 30:58]
  assign vertex_update_buffer_1_wr_en = apply_selecter_1_io_ddr_out_valid; // @[BFS.scala 294:40]
  assign vertex_update_buffer_1_rd_en = update_engine_1_io_xbar_in_ready; // @[BFS.scala 306:40]
  assign vertex_update_buffer_1_clk = clock; // @[BFS.scala 292:53]
  assign vertex_update_buffer_1_srst = reset; // @[BFS.scala 293:54]
  assign vertex_update_buffer_2_din = {apply_selecter_2_io_ddr_out_bits_tdata,io_level}; // @[Cat.scala 30:58]
  assign vertex_update_buffer_2_wr_en = apply_selecter_2_io_ddr_out_valid; // @[BFS.scala 294:40]
  assign vertex_update_buffer_2_rd_en = update_engine_2_io_xbar_in_ready; // @[BFS.scala 306:40]
  assign vertex_update_buffer_2_clk = clock; // @[BFS.scala 292:53]
  assign vertex_update_buffer_2_srst = reset; // @[BFS.scala 293:54]
  assign vertex_update_buffer_3_din = {apply_selecter_3_io_ddr_out_bits_tdata,io_level}; // @[Cat.scala 30:58]
  assign vertex_update_buffer_3_wr_en = apply_selecter_3_io_ddr_out_valid; // @[BFS.scala 294:40]
  assign vertex_update_buffer_3_rd_en = update_engine_3_io_xbar_in_ready; // @[BFS.scala 306:40]
  assign vertex_update_buffer_3_clk = clock; // @[BFS.scala 292:53]
  assign vertex_update_buffer_3_srst = reset; // @[BFS.scala 293:54]
  assign update_engine_0_clock = clock;
  assign update_engine_0_reset = reset;
  assign update_engine_0_io_axi_ddr_aw_ready = io_axi_0_ddr_aw_ready; // @[BFS.scala 305:17]
  assign update_engine_0_io_axi_ddr_w_ready = io_axi_0_ddr_w_ready; // @[BFS.scala 305:17]
  assign update_engine_0_io_xbar_in_valid = vertex_update_buffer_0_valid; // @[BFS.scala 301:41]
  assign update_engine_0_io_xbar_in_bits_tdata = vertex_update_buffer_0_dout[63:32]; // @[BFS.scala 298:80]
  assign update_engine_0_io_level_base_addr = io_level_base_addr; // @[BFS.scala 304:43]
  assign update_engine_0_io_level = vertex_update_buffer_0_dout[31:0]; // @[BFS.scala 302:67]
  assign update_engine_0_io_flush = io_flush & _update_engine_0_io_flush_T; // @[BFS.scala 303:45]
  assign update_engine_1_clock = clock;
  assign update_engine_1_reset = reset;
  assign update_engine_1_io_axi_ddr_aw_ready = io_axi_1_ddr_aw_ready; // @[BFS.scala 305:17]
  assign update_engine_1_io_axi_ddr_w_ready = io_axi_1_ddr_w_ready; // @[BFS.scala 305:17]
  assign update_engine_1_io_xbar_in_valid = vertex_update_buffer_1_valid; // @[BFS.scala 301:41]
  assign update_engine_1_io_xbar_in_bits_tdata = vertex_update_buffer_1_dout[63:32]; // @[BFS.scala 298:80]
  assign update_engine_1_io_level_base_addr = io_level_base_addr; // @[BFS.scala 304:43]
  assign update_engine_1_io_level = vertex_update_buffer_1_dout[31:0]; // @[BFS.scala 302:67]
  assign update_engine_1_io_flush = io_flush & _update_engine_1_io_flush_T; // @[BFS.scala 303:45]
  assign update_engine_2_clock = clock;
  assign update_engine_2_reset = reset;
  assign update_engine_2_io_axi_ddr_aw_ready = io_axi_2_ddr_aw_ready; // @[BFS.scala 305:17]
  assign update_engine_2_io_axi_ddr_w_ready = io_axi_2_ddr_w_ready; // @[BFS.scala 305:17]
  assign update_engine_2_io_xbar_in_valid = vertex_update_buffer_2_valid; // @[BFS.scala 301:41]
  assign update_engine_2_io_xbar_in_bits_tdata = vertex_update_buffer_2_dout[63:32]; // @[BFS.scala 298:80]
  assign update_engine_2_io_level_base_addr = io_level_base_addr; // @[BFS.scala 304:43]
  assign update_engine_2_io_level = vertex_update_buffer_2_dout[31:0]; // @[BFS.scala 302:67]
  assign update_engine_2_io_flush = io_flush & _update_engine_2_io_flush_T; // @[BFS.scala 303:45]
  assign update_engine_3_clock = clock;
  assign update_engine_3_reset = reset;
  assign update_engine_3_io_axi_ddr_aw_ready = io_axi_3_ddr_aw_ready; // @[BFS.scala 305:17]
  assign update_engine_3_io_axi_ddr_w_ready = io_axi_3_ddr_w_ready; // @[BFS.scala 305:17]
  assign update_engine_3_io_xbar_in_valid = vertex_update_buffer_3_valid; // @[BFS.scala 301:41]
  assign update_engine_3_io_xbar_in_bits_tdata = vertex_update_buffer_3_dout[63:32]; // @[BFS.scala 298:80]
  assign update_engine_3_io_level_base_addr = io_level_base_addr; // @[BFS.scala 304:43]
  assign update_engine_3_io_level = vertex_update_buffer_3_dout[31:0]; // @[BFS.scala 302:67]
  assign update_engine_3_io_flush = io_flush & _update_engine_3_io_flush_T; // @[BFS.scala 303:45]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 241:30]
      ready_counter <= 32'h0; // @[BFS.scala 241:30]
    end else if (~io_gather_in_ready & io_gather_in_valid) begin // @[BFS.scala 243:72]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 244:19]
    end
    if (reset) begin // @[BFS.scala 276:24]
      end_reg_0 <= 1'h0; // @[BFS.scala 276:24]
    end else begin
      end_reg_0 <= _GEN_1;
    end
    if (reset) begin // @[BFS.scala 276:24]
      end_reg_1 <= 1'h0; // @[BFS.scala 276:24]
    end else begin
      end_reg_1 <= _GEN_2;
    end
    if (reset) begin // @[BFS.scala 276:24]
      end_reg_2 <= 1'h0; // @[BFS.scala 276:24]
    end else begin
      end_reg_2 <= _GEN_3;
    end
    if (reset) begin // @[BFS.scala 276:24]
      end_reg_3 <= 1'h0; // @[BFS.scala 276:24]
    end else begin
      end_reg_3 <= _GEN_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ready_counter = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  end_reg_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  end_reg_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  end_reg_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  end_reg_3 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module regFile(
  input         clock,
  input         reset,
  input  [31:0] io_dataIn,
  output [31:0] io_dataOut,
  input         io_writeFlag,
  input  [4:0]  io_rptr,
  input  [4:0]  io_wptr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[util.scala 178:21]
  reg [31:0] regs_1; // @[util.scala 178:21]
  reg [31:0] regs_2; // @[util.scala 178:21]
  reg [31:0] regs_3; // @[util.scala 178:21]
  reg [31:0] regs_4; // @[util.scala 178:21]
  reg [31:0] regs_5; // @[util.scala 178:21]
  reg [31:0] regs_6; // @[util.scala 178:21]
  reg [31:0] regs_7; // @[util.scala 178:21]
  reg [31:0] regs_8; // @[util.scala 178:21]
  reg [31:0] regs_9; // @[util.scala 178:21]
  reg [31:0] regs_10; // @[util.scala 178:21]
  reg [31:0] regs_11; // @[util.scala 178:21]
  reg [31:0] regs_12; // @[util.scala 178:21]
  reg [31:0] regs_13; // @[util.scala 178:21]
  reg [31:0] regs_14; // @[util.scala 178:21]
  reg [31:0] regs_15; // @[util.scala 178:21]
  reg [31:0] regs_16; // @[util.scala 178:21]
  reg [31:0] regs_17; // @[util.scala 178:21]
  reg [31:0] regs_18; // @[util.scala 178:21]
  reg [31:0] regs_19; // @[util.scala 178:21]
  reg [31:0] regs_20; // @[util.scala 178:21]
  reg [31:0] regs_21; // @[util.scala 178:21]
  reg [31:0] regs_22; // @[util.scala 178:21]
  reg [31:0] regs_23; // @[util.scala 178:21]
  reg [31:0] regs_24; // @[util.scala 178:21]
  reg [31:0] regs_25; // @[util.scala 178:21]
  reg [31:0] regs_26; // @[util.scala 178:21]
  reg [31:0] regs_27; // @[util.scala 178:21]
  reg [31:0] regs_28; // @[util.scala 178:21]
  reg [31:0] regs_29; // @[util.scala 178:21]
  reg [31:0] regs_30; // @[util.scala 178:21]
  reg [31:0] regs_31; // @[util.scala 178:21]
  wire [31:0] _GEN_1 = 5'h1 == io_rptr ? regs_1 : regs_0; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_2 = 5'h2 == io_rptr ? regs_2 : _GEN_1; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_3 = 5'h3 == io_rptr ? regs_3 : _GEN_2; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_4 = 5'h4 == io_rptr ? regs_4 : _GEN_3; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_5 = 5'h5 == io_rptr ? regs_5 : _GEN_4; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_6 = 5'h6 == io_rptr ? regs_6 : _GEN_5; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_7 = 5'h7 == io_rptr ? regs_7 : _GEN_6; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_8 = 5'h8 == io_rptr ? regs_8 : _GEN_7; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_9 = 5'h9 == io_rptr ? regs_9 : _GEN_8; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_10 = 5'ha == io_rptr ? regs_10 : _GEN_9; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_11 = 5'hb == io_rptr ? regs_11 : _GEN_10; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_12 = 5'hc == io_rptr ? regs_12 : _GEN_11; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_13 = 5'hd == io_rptr ? regs_13 : _GEN_12; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_14 = 5'he == io_rptr ? regs_14 : _GEN_13; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_15 = 5'hf == io_rptr ? regs_15 : _GEN_14; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_16 = 5'h10 == io_rptr ? regs_16 : _GEN_15; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_17 = 5'h11 == io_rptr ? regs_17 : _GEN_16; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_18 = 5'h12 == io_rptr ? regs_18 : _GEN_17; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_19 = 5'h13 == io_rptr ? regs_19 : _GEN_18; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_20 = 5'h14 == io_rptr ? regs_20 : _GEN_19; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_21 = 5'h15 == io_rptr ? regs_21 : _GEN_20; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_22 = 5'h16 == io_rptr ? regs_22 : _GEN_21; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_23 = 5'h17 == io_rptr ? regs_23 : _GEN_22; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_24 = 5'h18 == io_rptr ? regs_24 : _GEN_23; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_25 = 5'h19 == io_rptr ? regs_25 : _GEN_24; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_26 = 5'h1a == io_rptr ? regs_26 : _GEN_25; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_27 = 5'h1b == io_rptr ? regs_27 : _GEN_26; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_28 = 5'h1c == io_rptr ? regs_28 : _GEN_27; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_29 = 5'h1d == io_rptr ? regs_29 : _GEN_28; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_30 = 5'h1e == io_rptr ? regs_30 : _GEN_29; // @[util.scala 180:14 util.scala 180:14]
  assign io_dataOut = 5'h1f == io_rptr ? regs_31 : _GEN_30; // @[util.scala 180:14 util.scala 180:14]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 178:21]
      regs_0 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h0 == io_wptr) begin // @[util.scala 183:19]
        regs_0 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_1 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1 == io_wptr) begin // @[util.scala 183:19]
        regs_1 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_2 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h2 == io_wptr) begin // @[util.scala 183:19]
        regs_2 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_3 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h3 == io_wptr) begin // @[util.scala 183:19]
        regs_3 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_4 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h4 == io_wptr) begin // @[util.scala 183:19]
        regs_4 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_5 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h5 == io_wptr) begin // @[util.scala 183:19]
        regs_5 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_6 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h6 == io_wptr) begin // @[util.scala 183:19]
        regs_6 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_7 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h7 == io_wptr) begin // @[util.scala 183:19]
        regs_7 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_8 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h8 == io_wptr) begin // @[util.scala 183:19]
        regs_8 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_9 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h9 == io_wptr) begin // @[util.scala 183:19]
        regs_9 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_10 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'ha == io_wptr) begin // @[util.scala 183:19]
        regs_10 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_11 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hb == io_wptr) begin // @[util.scala 183:19]
        regs_11 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_12 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hc == io_wptr) begin // @[util.scala 183:19]
        regs_12 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_13 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hd == io_wptr) begin // @[util.scala 183:19]
        regs_13 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_14 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'he == io_wptr) begin // @[util.scala 183:19]
        regs_14 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_15 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hf == io_wptr) begin // @[util.scala 183:19]
        regs_15 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_16 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h10 == io_wptr) begin // @[util.scala 183:19]
        regs_16 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_17 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h11 == io_wptr) begin // @[util.scala 183:19]
        regs_17 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_18 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h12 == io_wptr) begin // @[util.scala 183:19]
        regs_18 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_19 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h13 == io_wptr) begin // @[util.scala 183:19]
        regs_19 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_20 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h14 == io_wptr) begin // @[util.scala 183:19]
        regs_20 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_21 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h15 == io_wptr) begin // @[util.scala 183:19]
        regs_21 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_22 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h16 == io_wptr) begin // @[util.scala 183:19]
        regs_22 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_23 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h17 == io_wptr) begin // @[util.scala 183:19]
        regs_23 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_24 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h18 == io_wptr) begin // @[util.scala 183:19]
        regs_24 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_25 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h19 == io_wptr) begin // @[util.scala 183:19]
        regs_25 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_26 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1a == io_wptr) begin // @[util.scala 183:19]
        regs_26 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_27 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1b == io_wptr) begin // @[util.scala 183:19]
        regs_27 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_28 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1c == io_wptr) begin // @[util.scala 183:19]
        regs_28 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_29 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1d == io_wptr) begin // @[util.scala 183:19]
        regs_29 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_30 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1e == io_wptr) begin // @[util.scala 183:19]
        regs_30 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_31 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1f == io_wptr) begin // @[util.scala 183:19]
        regs_31 <= io_dataIn; // @[util.scala 183:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module regFile_1(
  input         clock,
  input         reset,
  input  [63:0] io_dataIn,
  output [63:0] io_dataOut,
  input         io_writeFlag,
  input  [4:0]  io_rptr,
  input  [4:0]  io_wptr
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0; // @[util.scala 178:21]
  reg [63:0] regs_1; // @[util.scala 178:21]
  reg [63:0] regs_2; // @[util.scala 178:21]
  reg [63:0] regs_3; // @[util.scala 178:21]
  reg [63:0] regs_4; // @[util.scala 178:21]
  reg [63:0] regs_5; // @[util.scala 178:21]
  reg [63:0] regs_6; // @[util.scala 178:21]
  reg [63:0] regs_7; // @[util.scala 178:21]
  reg [63:0] regs_8; // @[util.scala 178:21]
  reg [63:0] regs_9; // @[util.scala 178:21]
  reg [63:0] regs_10; // @[util.scala 178:21]
  reg [63:0] regs_11; // @[util.scala 178:21]
  reg [63:0] regs_12; // @[util.scala 178:21]
  reg [63:0] regs_13; // @[util.scala 178:21]
  reg [63:0] regs_14; // @[util.scala 178:21]
  reg [63:0] regs_15; // @[util.scala 178:21]
  reg [63:0] regs_16; // @[util.scala 178:21]
  reg [63:0] regs_17; // @[util.scala 178:21]
  reg [63:0] regs_18; // @[util.scala 178:21]
  reg [63:0] regs_19; // @[util.scala 178:21]
  reg [63:0] regs_20; // @[util.scala 178:21]
  reg [63:0] regs_21; // @[util.scala 178:21]
  reg [63:0] regs_22; // @[util.scala 178:21]
  reg [63:0] regs_23; // @[util.scala 178:21]
  reg [63:0] regs_24; // @[util.scala 178:21]
  reg [63:0] regs_25; // @[util.scala 178:21]
  reg [63:0] regs_26; // @[util.scala 178:21]
  reg [63:0] regs_27; // @[util.scala 178:21]
  reg [63:0] regs_28; // @[util.scala 178:21]
  reg [63:0] regs_29; // @[util.scala 178:21]
  reg [63:0] regs_30; // @[util.scala 178:21]
  reg [63:0] regs_31; // @[util.scala 178:21]
  wire [63:0] _GEN_1 = 5'h1 == io_rptr ? regs_1 : regs_0; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_2 = 5'h2 == io_rptr ? regs_2 : _GEN_1; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_3 = 5'h3 == io_rptr ? regs_3 : _GEN_2; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_4 = 5'h4 == io_rptr ? regs_4 : _GEN_3; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_5 = 5'h5 == io_rptr ? regs_5 : _GEN_4; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_6 = 5'h6 == io_rptr ? regs_6 : _GEN_5; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_7 = 5'h7 == io_rptr ? regs_7 : _GEN_6; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_8 = 5'h8 == io_rptr ? regs_8 : _GEN_7; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_9 = 5'h9 == io_rptr ? regs_9 : _GEN_8; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_10 = 5'ha == io_rptr ? regs_10 : _GEN_9; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_11 = 5'hb == io_rptr ? regs_11 : _GEN_10; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_12 = 5'hc == io_rptr ? regs_12 : _GEN_11; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_13 = 5'hd == io_rptr ? regs_13 : _GEN_12; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_14 = 5'he == io_rptr ? regs_14 : _GEN_13; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_15 = 5'hf == io_rptr ? regs_15 : _GEN_14; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_16 = 5'h10 == io_rptr ? regs_16 : _GEN_15; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_17 = 5'h11 == io_rptr ? regs_17 : _GEN_16; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_18 = 5'h12 == io_rptr ? regs_18 : _GEN_17; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_19 = 5'h13 == io_rptr ? regs_19 : _GEN_18; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_20 = 5'h14 == io_rptr ? regs_20 : _GEN_19; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_21 = 5'h15 == io_rptr ? regs_21 : _GEN_20; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_22 = 5'h16 == io_rptr ? regs_22 : _GEN_21; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_23 = 5'h17 == io_rptr ? regs_23 : _GEN_22; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_24 = 5'h18 == io_rptr ? regs_24 : _GEN_23; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_25 = 5'h19 == io_rptr ? regs_25 : _GEN_24; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_26 = 5'h1a == io_rptr ? regs_26 : _GEN_25; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_27 = 5'h1b == io_rptr ? regs_27 : _GEN_26; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_28 = 5'h1c == io_rptr ? regs_28 : _GEN_27; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_29 = 5'h1d == io_rptr ? regs_29 : _GEN_28; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_30 = 5'h1e == io_rptr ? regs_30 : _GEN_29; // @[util.scala 180:14 util.scala 180:14]
  assign io_dataOut = 5'h1f == io_rptr ? regs_31 : _GEN_30; // @[util.scala 180:14 util.scala 180:14]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 178:21]
      regs_0 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h0 == io_wptr) begin // @[util.scala 183:19]
        regs_0 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_1 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1 == io_wptr) begin // @[util.scala 183:19]
        regs_1 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_2 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h2 == io_wptr) begin // @[util.scala 183:19]
        regs_2 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_3 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h3 == io_wptr) begin // @[util.scala 183:19]
        regs_3 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_4 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h4 == io_wptr) begin // @[util.scala 183:19]
        regs_4 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_5 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h5 == io_wptr) begin // @[util.scala 183:19]
        regs_5 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_6 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h6 == io_wptr) begin // @[util.scala 183:19]
        regs_6 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_7 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h7 == io_wptr) begin // @[util.scala 183:19]
        regs_7 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_8 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h8 == io_wptr) begin // @[util.scala 183:19]
        regs_8 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_9 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h9 == io_wptr) begin // @[util.scala 183:19]
        regs_9 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_10 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'ha == io_wptr) begin // @[util.scala 183:19]
        regs_10 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_11 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hb == io_wptr) begin // @[util.scala 183:19]
        regs_11 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_12 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hc == io_wptr) begin // @[util.scala 183:19]
        regs_12 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_13 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hd == io_wptr) begin // @[util.scala 183:19]
        regs_13 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_14 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'he == io_wptr) begin // @[util.scala 183:19]
        regs_14 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_15 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hf == io_wptr) begin // @[util.scala 183:19]
        regs_15 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_16 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h10 == io_wptr) begin // @[util.scala 183:19]
        regs_16 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_17 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h11 == io_wptr) begin // @[util.scala 183:19]
        regs_17 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_18 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h12 == io_wptr) begin // @[util.scala 183:19]
        regs_18 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_19 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h13 == io_wptr) begin // @[util.scala 183:19]
        regs_19 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_20 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h14 == io_wptr) begin // @[util.scala 183:19]
        regs_20 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_21 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h15 == io_wptr) begin // @[util.scala 183:19]
        regs_21 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_22 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h16 == io_wptr) begin // @[util.scala 183:19]
        regs_22 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_23 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h17 == io_wptr) begin // @[util.scala 183:19]
        regs_23 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_24 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h18 == io_wptr) begin // @[util.scala 183:19]
        regs_24 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_25 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h19 == io_wptr) begin // @[util.scala 183:19]
        regs_25 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_26 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1a == io_wptr) begin // @[util.scala 183:19]
        regs_26 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_27 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1b == io_wptr) begin // @[util.scala 183:19]
        regs_27 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_28 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1c == io_wptr) begin // @[util.scala 183:19]
        regs_28 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_29 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1d == io_wptr) begin // @[util.scala 183:19]
        regs_29 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_30 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1e == io_wptr) begin // @[util.scala 183:19]
        regs_30 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_31 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1f == io_wptr) begin // @[util.scala 183:19]
        regs_31 <= io_dataIn; // @[util.scala 183:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regs_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regs_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regs_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regs_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regs_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regs_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regs_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regs_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regs_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regs_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regs_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regs_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regs_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regs_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regs_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regs_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regs_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regs_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regs_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regs_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regs_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regs_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regs_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regs_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regs_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regs_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regs_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regs_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regs_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regs_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module readEdge_engine(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_rdata,
  input  [5:0]   io_in_bits_rid,
  input          io_in_bits_rlast,
  input          io_out_ready,
  output         io_out_valid,
  output [63:0]  io_out_bits_araddr,
  output [5:0]   io_out_bits_arid,
  output [7:0]   io_out_bits_arlen,
  output [2:0]   io_out_bits_arsize,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_edge_base_addr,
  output         io_read_edge_fifo_empty,
  output [7:0]   io_credit,
  input          io_credit_req_valid,
  input  [5:0]   io_credit_req_bits_arid,
  input  [31:0]  io_credit_req_bits_vid,
  output [63:0]  io_traveled_edges,
  input          io_signal
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  rid2vid_clock; // @[BFS.scala 468:23]
  wire  rid2vid_reset; // @[BFS.scala 468:23]
  wire [31:0] rid2vid_io_dataIn; // @[BFS.scala 468:23]
  wire [31:0] rid2vid_io_dataOut; // @[BFS.scala 468:23]
  wire  rid2vid_io_writeFlag; // @[BFS.scala 468:23]
  wire [4:0] rid2vid_io_rptr; // @[BFS.scala 468:23]
  wire [4:0] rid2vid_io_wptr; // @[BFS.scala 468:23]
  wire  num_regfile_clock; // @[BFS.scala 474:27]
  wire  num_regfile_reset; // @[BFS.scala 474:27]
  wire [63:0] num_regfile_io_dataIn; // @[BFS.scala 474:27]
  wire [63:0] num_regfile_io_dataOut; // @[BFS.scala 474:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 474:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 474:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 474:27]
  wire  edge_read_buffer__full; // @[BFS.scala 524:32]
  wire [71:0] edge_read_buffer__din; // @[BFS.scala 524:32]
  wire  edge_read_buffer__wr_en; // @[BFS.scala 524:32]
  wire  edge_read_buffer__empty; // @[BFS.scala 524:32]
  wire [71:0] edge_read_buffer__dout; // @[BFS.scala 524:32]
  wire  edge_read_buffer__rd_en; // @[BFS.scala 524:32]
  wire [5:0] edge_read_buffer__data_count; // @[BFS.scala 524:32]
  wire  edge_read_buffer__clk; // @[BFS.scala 524:32]
  wire  edge_read_buffer__srst; // @[BFS.scala 524:32]
  wire  edge_read_buffer__valid; // @[BFS.scala 524:32]
  wire  free_queue_full; // @[BFS.scala 574:26]
  wire [5:0] free_queue_din; // @[BFS.scala 574:26]
  wire  free_queue_wr_en; // @[BFS.scala 574:26]
  wire  free_queue_empty; // @[BFS.scala 574:26]
  wire [5:0] free_queue_dout; // @[BFS.scala 574:26]
  wire  free_queue_rd_en; // @[BFS.scala 574:26]
  wire [5:0] free_queue_data_count; // @[BFS.scala 574:26]
  wire  free_queue_clk; // @[BFS.scala 574:26]
  wire  free_queue_srst; // @[BFS.scala 574:26]
  wire  free_queue_valid; // @[BFS.scala 574:26]
  reg [1:0] status; // @[BFS.scala 445:23]
  wire  _T = status == 2'h0; // @[BFS.scala 446:15]
  wire  _T_2 = status == 2'h0 & io_in_valid & io_in_ready; // @[BFS.scala 446:48]
  wire  _T_6 = status == 2'h2; // @[BFS.scala 454:22]
  wire  _T_7 = status == 2'h1; // @[BFS.scala 454:60]
  wire  _T_8 = status == 2'h2 | status == 2'h1; // @[BFS.scala 454:50]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 458:35]
  wire  _T_13 = io_in_valid & io_in_ready; // @[BFS.scala 461:26]
  wire  _T_16 = ~io_in_bits_rid[5]; // @[BFS.scala 461:44]
  wire  _T_17 = io_in_valid & io_in_ready & ~io_in_bits_rid[5]; // @[BFS.scala 461:41]
  wire [63:0] _GEN_131 = {{32'd0}, io_in_bits_rdata[63:32]}; // @[BFS.scala 463:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_131; // @[BFS.scala 463:46]
  reg [31:0] num; // @[BFS.scala 475:20]
  wire [31:0] _num_T_4 = num_regfile_io_dataOut[63:32] - 32'h4; // @[BFS.scala 479:103]
  wire [31:0] _num_T_10 = io_in_bits_rdata[63:32] - 32'h2; // @[BFS.scala 482:42]
  wire [31:0] _num_T_13 = num - 32'h4; // @[BFS.scala 488:18]
  wire [31:0] _num_T_17 = num > 32'h4 ? _num_T_13 : 32'h0; // @[BFS.scala 494:17]
  wire [31:0] _GEN_8 = io_in_bits_rlast ? 32'h0 : _num_T_17; // @[BFS.scala 491:36 BFS.scala 492:11 BFS.scala 494:11]
  wire  _T_44 = _T & _T_16; // @[BFS.scala 504:43]
  wire  _GEN_12 = _T_8 & num > 32'h0; // @[BFS.scala 510:94 BFS.scala 511:11 BFS.scala 501:9]
  wire  _GEN_13 = _T & _T_16 ? 1'h0 : _GEN_12; // @[BFS.scala 504:72 BFS.scala 506:13]
  wire  keep_0 = _T & io_in_bits_rid[5] ? num_regfile_io_dataOut[63:32] > 32'h0 : _GEN_13; // @[BFS.scala 502:65 BFS.scala 503:11]
  wire  _GEN_15 = _T_8 & num > 32'h1; // @[BFS.scala 510:94 BFS.scala 511:11 BFS.scala 501:9]
  wire  _GEN_16 = _T & _T_16 ? 1'h0 : _GEN_15; // @[BFS.scala 504:72 BFS.scala 506:13]
  wire  keep_1 = _T & io_in_bits_rid[5] ? num_regfile_io_dataOut[63:32] > 32'h1 : _GEN_16; // @[BFS.scala 502:65 BFS.scala 503:11]
  wire  _GEN_18 = _T_8 & num > 32'h2; // @[BFS.scala 510:94 BFS.scala 511:11 BFS.scala 501:9]
  wire  _GEN_19 = _T & _T_16 ? io_in_bits_rdata[63:32] > 32'h0 : _GEN_18; // @[BFS.scala 504:72 BFS.scala 508:13]
  wire  keep_2 = _T & io_in_bits_rid[5] ? num_regfile_io_dataOut[63:32] > 32'h2 : _GEN_19; // @[BFS.scala 502:65 BFS.scala 503:11]
  wire  _GEN_21 = _T_8 & num > 32'h3; // @[BFS.scala 510:94 BFS.scala 511:11 BFS.scala 501:9]
  wire  _GEN_22 = _T & _T_16 ? io_in_bits_rdata[63:32] > 32'h1 : _GEN_21; // @[BFS.scala 504:72 BFS.scala 508:13]
  wire  keep_3 = _T & io_in_bits_rid[5] ? num_regfile_io_dataOut[63:32] > 32'h3 : _GEN_22; // @[BFS.scala 502:65 BFS.scala 503:11]
  wire [95:0] io_xbar_out_bits_tdata_hi = io_in_bits_rdata[127:32]; // @[BFS.scala 518:51]
  wire [127:0] _io_xbar_out_bits_tdata_T = {io_xbar_out_bits_tdata_hi,rid2vid_io_dataOut}; // @[Cat.scala 30:58]
  wire [1:0] io_xbar_out_bits_tkeep_lo = {keep_1,keep_0}; // @[BFS.scala 521:40]
  wire [1:0] io_xbar_out_bits_tkeep_hi = {keep_3,keep_2}; // @[BFS.scala 521:40]
  wire [31:0] _edge_read_buffer_din_count_T_3 = io_in_bits_rdata[63:32] - 32'he; // @[BFS.scala 529:73]
  wire [31:0] _edge_read_buffer_din_index_T_4 = num_regfile_io_dataOut[31:0] + 32'h40; // @[BFS.scala 545:56]
  wire [31:0] _GEN_26 = num_regfile_io_dataOut[63:32] > 32'h40 ? _edge_read_buffer_din_index_T_4 : io_in_bits_rdata[31:0
    ]; // @[BFS.scala 541:85 BFS.scala 544:36 BFS.scala 530:30]
  wire [31:0] _GEN_31 = io_in_bits_rid[5] ? _GEN_26 : io_in_bits_rdata[31:0]; // @[BFS.scala 538:35 BFS.scala 530:30]
  wire [31:0] edge_read_buffer_din_index = _T_13 & _T ? _GEN_31 : io_in_bits_rdata[31:0]; // @[BFS.scala 536:64 BFS.scala 530:30]
  wire [4:0] _GEN_29 = io_in_bits_rid[5] ? io_in_bits_rid[4:0] : 5'h0; // @[BFS.scala 538:35 BFS.scala 540:36 BFS.scala 532:32]
  wire [4:0] _GEN_34 = _T_13 & _T ? _GEN_29 : 5'h0; // @[BFS.scala 536:64 BFS.scala 532:32]
  wire [5:0] edge_read_buffer_din_reg_ptr = {{1'd0}, _GEN_34}; // @[BFS.scala 526:34]
  wire [31:0] _edge_read_buffer_din_count_T_6 = num_regfile_io_dataOut[63:32] - 32'h40; // @[BFS.scala 543:50]
  wire [31:0] _GEN_25 = num_regfile_io_dataOut[63:32] > 32'h40 ? _edge_read_buffer_din_count_T_6 : 32'h0; // @[BFS.scala 541:85 BFS.scala 542:36 BFS.scala 547:36]
  wire [31:0] _GEN_27 = io_in_bits_rdata[63:32] < 32'he ? 32'h0 : _edge_read_buffer_din_count_T_3; // @[BFS.scala 550:66 BFS.scala 551:36 BFS.scala 529:30]
  wire [31:0] _GEN_30 = io_in_bits_rid[5] ? _GEN_25 : _GEN_27; // @[BFS.scala 538:35]
  wire [31:0] edge_read_buffer_din_count = _T_13 & _T ? _GEN_30 : _edge_read_buffer_din_count_T_3; // @[BFS.scala 536:64 BFS.scala 529:30]
  wire  _GEN_28 = io_in_bits_rid[5] ? 1'h0 : 1'h1; // @[BFS.scala 538:35 BFS.scala 539:35 BFS.scala 531:31]
  wire  edge_read_buffer_din_is_new = _T_13 & _T ? _GEN_28 : 1'h1; // @[BFS.scala 536:64 BFS.scala 531:31]
  wire [70:0] _edge_read_buffer_io_din_T = {edge_read_buffer_din_count,edge_read_buffer_din_is_new,
    edge_read_buffer_din_index,edge_read_buffer_din_reg_ptr}; // @[BFS.scala 535:57]
  wire [5:0] edge_read_buffer_dout_reg_ptr = edge_read_buffer__dout[5:0]; // @[BFS.scala 558:65]
  wire [31:0] edge_read_buffer_dout_index = edge_read_buffer__dout[37:6]; // @[BFS.scala 558:65]
  wire  edge_read_buffer_dout_is_new = edge_read_buffer__dout[38]; // @[BFS.scala 558:65]
  wire [31:0] edge_read_buffer_dout_count = edge_read_buffer__dout[70:39]; // @[BFS.scala 558:65]
  reg [3:0] cache_status; // @[BFS.scala 573:29]
  reg [5:0] init_seq; // @[BFS.scala 575:25]
  wire  _T_98 = cache_status == 4'h6; // @[BFS.scala 576:21]
  wire [5:0] _init_seq_T_1 = init_seq + 6'h1; // @[BFS.scala 577:26]
  reg [31:0] expand_index; // @[BFS.scala 579:29]
  reg [31:0] expand_count; // @[BFS.scala 580:29]
  reg [31:0] credit; // @[BFS.scala 581:23]
  wire  _T_105 = cache_status == 4'h0; // @[BFS.scala 586:27]
  wire  _T_108 = edge_read_buffer_dout_count == 32'h0; // @[BFS.scala 588:29]
  wire  _T_111 = edge_read_buffer_dout_count > 32'h40 & credit > 32'h4; // @[BFS.scala 591:65]
  wire [2:0] _GEN_38 = edge_read_buffer_dout_count > 32'h40 & credit > 32'h4 ? 3'h5 : 3'h2; // @[BFS.scala 591:99 BFS.scala 592:24 BFS.scala 596:24]
  wire [31:0] _GEN_39 = edge_read_buffer_dout_count > 32'h40 & credit > 32'h4 ? edge_read_buffer_dout_index :
    expand_index; // @[BFS.scala 591:99 BFS.scala 593:24 BFS.scala 579:29]
  wire [31:0] _GEN_40 = edge_read_buffer_dout_count > 32'h40 & credit > 32'h4 ? edge_read_buffer_dout_count :
    expand_count; // @[BFS.scala 591:99 BFS.scala 594:24 BFS.scala 580:29]
  wire [2:0] _GEN_41 = edge_read_buffer_dout_count == 32'h0 ? 3'h7 : _GEN_38; // @[BFS.scala 588:37 BFS.scala 589:22]
  wire [31:0] _GEN_42 = edge_read_buffer_dout_count == 32'h0 ? expand_index : _GEN_39; // @[BFS.scala 588:37 BFS.scala 579:29]
  wire [31:0] _GEN_43 = edge_read_buffer_dout_count == 32'h0 ? expand_count : _GEN_40; // @[BFS.scala 588:37 BFS.scala 580:29]
  wire [1:0] _GEN_44 = _T_111 ? 2'h1 : 2'h3; // @[BFS.scala 603:99 BFS.scala 604:24 BFS.scala 608:24]
  wire [2:0] _GEN_47 = _T_108 ? 3'h4 : {{1'd0}, _GEN_44}; // @[BFS.scala 600:37 BFS.scala 601:22]
  wire [2:0] _GEN_50 = edge_read_buffer_dout_is_new ? _GEN_41 : _GEN_47; // @[BFS.scala 587:50]
  wire [31:0] _GEN_51 = edge_read_buffer_dout_is_new ? _GEN_42 : _GEN_42; // @[BFS.scala 587:50]
  wire [31:0] _GEN_52 = edge_read_buffer_dout_is_new ? _GEN_43 : _GEN_43; // @[BFS.scala 587:50]
  wire  _T_116 = io_out_ready & io_out_valid; // @[BFS.scala 612:27]
  wire  _T_117 = cache_status == 4'h2; // @[BFS.scala 612:59]
  wire  _T_120 = cache_status == 4'h3; // @[BFS.scala 615:59]
  wire  _T_122 = cache_status == 4'h7; // @[BFS.scala 618:27]
  wire  _T_123 = cache_status == 4'h4; // @[BFS.scala 621:27]
  wire  _T_125 = cache_status == 4'h5; // @[BFS.scala 624:59]
  wire  _T_126 = _T_116 & cache_status == 4'h5; // @[BFS.scala 624:43]
  wire [31:0] _expand_index_T_1 = expand_index + 32'h40; // @[BFS.scala 625:34]
  wire [31:0] _expand_count_T_1 = expand_count - 32'h40; // @[BFS.scala 626:34]
  wire  _T_130 = credit <= 32'h4 | expand_count <= 32'h80; // @[BFS.scala 627:42]
  wire [3:0] _GEN_53 = credit <= 32'h4 | expand_count <= 32'h80 ? 4'h8 : cache_status; // @[BFS.scala 627:111 BFS.scala 628:20 BFS.scala 573:29]
  wire  _T_132 = cache_status == 4'h1; // @[BFS.scala 630:59]
  wire  _T_133 = _T_116 & cache_status == 4'h1; // @[BFS.scala 630:43]
  wire [3:0] _GEN_54 = _T_130 ? 4'h8 : 4'h5; // @[BFS.scala 633:111 BFS.scala 634:20 BFS.scala 636:20]
  wire  _T_139 = cache_status == 4'h8; // @[BFS.scala 638:59]
  wire  _T_140 = _T_116 & cache_status == 4'h8; // @[BFS.scala 638:43]
  wire [3:0] _GEN_55 = _T_116 & cache_status == 4'h8 ? 4'h0 : cache_status; // @[BFS.scala 638:83 BFS.scala 639:18 BFS.scala 573:29]
  wire [31:0] _GEN_57 = _T_116 & cache_status == 4'h1 ? _expand_index_T_1 : expand_index; // @[BFS.scala 630:91 BFS.scala 631:18 BFS.scala 579:29]
  wire [31:0] _GEN_58 = _T_116 & cache_status == 4'h1 ? _expand_count_T_1 : expand_count; // @[BFS.scala 630:91 BFS.scala 632:18 BFS.scala 580:29]
  wire [3:0] _GEN_59 = _T_116 & cache_status == 4'h1 ? _GEN_54 : _GEN_55; // @[BFS.scala 630:91]
  wire  _GEN_60 = _T_116 & cache_status == 4'h1 ? 1'h0 : _T_140; // @[BFS.scala 630:91 BFS.scala 534:29]
  wire [31:0] _GEN_61 = _T_116 & cache_status == 4'h5 ? _expand_index_T_1 : _GEN_57; // @[BFS.scala 624:91 BFS.scala 625:18]
  wire [31:0] _GEN_62 = _T_116 & cache_status == 4'h5 ? _expand_count_T_1 : _GEN_58; // @[BFS.scala 624:91 BFS.scala 626:18]
  wire [3:0] _GEN_63 = _T_116 & cache_status == 4'h5 ? _GEN_53 : _GEN_59; // @[BFS.scala 624:91]
  wire  _GEN_64 = _T_116 & cache_status == 4'h5 ? 1'h0 : _GEN_60; // @[BFS.scala 624:91 BFS.scala 534:29]
  wire [3:0] _GEN_65 = cache_status == 4'h4 ? 4'h0 : _GEN_63; // @[BFS.scala 621:51 BFS.scala 622:18]
  wire  _GEN_66 = cache_status == 4'h4 | _GEN_64; // @[BFS.scala 621:51 BFS.scala 623:31]
  wire [31:0] _GEN_67 = cache_status == 4'h4 ? expand_index : _GEN_61; // @[BFS.scala 621:51 BFS.scala 579:29]
  wire [31:0] _GEN_68 = cache_status == 4'h4 ? expand_count : _GEN_62; // @[BFS.scala 621:51 BFS.scala 580:29]
  wire [3:0] _GEN_69 = cache_status == 4'h7 ? 4'h0 : _GEN_65; // @[BFS.scala 618:55 BFS.scala 619:18]
  wire  _GEN_70 = cache_status == 4'h7 | _GEN_66; // @[BFS.scala 618:55 BFS.scala 620:31]
  wire [31:0] _GEN_71 = cache_status == 4'h7 ? expand_index : _GEN_67; // @[BFS.scala 618:55 BFS.scala 579:29]
  wire [31:0] _GEN_72 = cache_status == 4'h7 ? expand_count : _GEN_68; // @[BFS.scala 618:55 BFS.scala 580:29]
  wire [3:0] _GEN_73 = _T_116 & cache_status == 4'h3 ? 4'h0 : _GEN_69; // @[BFS.scala 615:87 BFS.scala 616:18]
  wire  _GEN_74 = _T_116 & cache_status == 4'h3 | _GEN_70; // @[BFS.scala 615:87 BFS.scala 617:31]
  wire [31:0] _GEN_75 = _T_116 & cache_status == 4'h3 ? expand_index : _GEN_71; // @[BFS.scala 615:87 BFS.scala 579:29]
  wire [31:0] _GEN_76 = _T_116 & cache_status == 4'h3 ? expand_count : _GEN_72; // @[BFS.scala 615:87 BFS.scala 580:29]
  wire [3:0] _GEN_77 = io_out_ready & io_out_valid & cache_status == 4'h2 ? 4'h0 : _GEN_73; // @[BFS.scala 612:84 BFS.scala 613:18]
  wire  _GEN_78 = io_out_ready & io_out_valid & cache_status == 4'h2 | _GEN_74; // @[BFS.scala 612:84 BFS.scala 614:31]
  wire [31:0] _GEN_79 = io_out_ready & io_out_valid & cache_status == 4'h2 ? expand_index : _GEN_75; // @[BFS.scala 612:84 BFS.scala 579:29]
  wire [31:0] _GEN_80 = io_out_ready & io_out_valid & cache_status == 4'h2 ? expand_count : _GEN_76; // @[BFS.scala 612:84 BFS.scala 580:29]
  wire  _GEN_84 = cache_status == 4'h0 & edge_read_buffer__valid ? 1'h0 : _GEN_78; // @[BFS.scala 586:77 BFS.scala 534:29]
  wire  _GEN_88 = _T_98 & init_seq == 6'h1f ? 1'h0 : _GEN_84; // @[BFS.scala 584:77 BFS.scala 534:29]
  wire  _num_vertex_T_2 = _T_139 & expand_count <= 32'h40; // @[BFS.scala 645:43]
  wire  _num_vertex_T_3 = edge_read_buffer_dout_count <= 32'h40; // @[BFS.scala 647:23]
  wire [31:0] _num_vertex_T_4 = _num_vertex_T_3 ? edge_read_buffer_dout_count : 32'h40; // @[Mux.scala 98:16]
  wire [31:0] num_vertex = _num_vertex_T_2 ? expand_count : _num_vertex_T_4; // @[Mux.scala 98:16]
  wire [31:0] _arlen_T_1 = {num_vertex[31:2], 2'h0}; // @[BFS.scala 649:63]
  wire [29:0] _arlen_T_6 = num_vertex[31:2] - 30'h1; // @[BFS.scala 651:57]
  wire [29:0] arlen = _arlen_T_1 < num_vertex ? num_vertex[31:2] : _arlen_T_6; // @[BFS.scala 649:18]
  wire [31:0] _io_out_bits_araddr_T_5 = _T_139 | _T_125 | _T_132 ? expand_index : edge_read_buffer_dout_index; // @[BFS.scala 654:11]
  wire [33:0] _GEN_132 = {_io_out_bits_araddr_T_5, 2'h0}; // @[BFS.scala 656:52]
  wire [34:0] _io_out_bits_araddr_T_6 = {{1'd0}, _GEN_132}; // @[BFS.scala 656:52]
  wire [63:0] _GEN_133 = {{29'd0}, _io_out_bits_araddr_T_6}; // @[BFS.scala 653:23]
  wire  _io_out_valid_T_4 = _T_117 | _T_120 | _T_139; // @[BFS.scala 657:100]
  wire  _io_out_bits_arsize_T = num_vertex <= 32'h1; // @[BFS.scala 664:23]
  wire  _io_out_bits_arsize_T_1 = num_vertex <= 32'h2; // @[BFS.scala 664:23]
  wire [2:0] _io_out_bits_arsize_T_2 = _io_out_bits_arsize_T_1 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  wire [4:0] io_out_bits_arid_lo = _T_117 | _T_125 | _T_139 ? free_queue_dout[4:0] : edge_read_buffer_dout_reg_ptr[4:0]; // @[BFS.scala 667:8]
  wire  _num_regfile_io_writeFlag_T_1 = free_queue_valid & io_out_ready & io_out_valid; // @[BFS.scala 684:71]
  wire [63:0] _num_regfile_io_dataIn_T = {edge_read_buffer_dout_count,edge_read_buffer_dout_index}; // @[Cat.scala 30:58]
  wire [38:0] _num_regfile_io_dataIn_T_2 = {7'h40,expand_index}; // @[Cat.scala 30:58]
  wire [63:0] _num_regfile_io_dataIn_T_4 = {expand_count,expand_index}; // @[Cat.scala 30:58]
  wire [5:0] _GEN_93 = _T_139 ? free_queue_dout : 6'h0; // @[BFS.scala 709:51 BFS.scala 710:25 BFS.scala 673:23]
  wire  _GEN_94 = _T_139 & _T_116; // @[BFS.scala 709:51 BFS.scala 711:25 BFS.scala 678:23]
  wire  _GEN_95 = _T_139 & _num_regfile_io_writeFlag_T_1; // @[BFS.scala 709:51 BFS.scala 712:30 BFS.scala 672:28]
  wire [63:0] _GEN_96 = _T_139 ? _num_regfile_io_dataIn_T_4 : 64'h0; // @[BFS.scala 709:51 BFS.scala 713:27 BFS.scala 674:25]
  wire [5:0] _GEN_97 = _T_132 ? edge_read_buffer_dout_reg_ptr : _GEN_93; // @[BFS.scala 704:59 BFS.scala 705:25]
  wire  _GEN_98 = _T_132 ? _T_116 : _GEN_95; // @[BFS.scala 704:59 BFS.scala 706:30]
  wire [63:0] _GEN_99 = _T_132 ? {{25'd0}, _num_regfile_io_dataIn_T_2} : _GEN_96; // @[BFS.scala 704:59 BFS.scala 707:27]
  wire  _GEN_100 = _T_132 ? 1'h0 : _GEN_94; // @[BFS.scala 704:59 BFS.scala 678:23]
  wire [5:0] _GEN_101 = _T_125 ? free_queue_dout : _GEN_97; // @[BFS.scala 698:59 BFS.scala 699:25]
  wire  _GEN_102 = _T_125 ? _T_116 : _GEN_100; // @[BFS.scala 698:59 BFS.scala 700:25]
  wire  _GEN_103 = _T_125 ? _num_regfile_io_writeFlag_T_1 : _GEN_98; // @[BFS.scala 698:59 BFS.scala 701:30]
  wire [63:0] _GEN_104 = _T_125 ? {{25'd0}, _num_regfile_io_dataIn_T_2} : _GEN_99; // @[BFS.scala 698:59 BFS.scala 702:27]
  wire [5:0] _GEN_105 = _T_98 ? init_seq : 6'h0; // @[BFS.scala 695:56 BFS.scala 696:23 BFS.scala 679:21]
  wire [5:0] _GEN_107 = _T_98 ? 6'h0 : _GEN_101; // @[BFS.scala 695:56 BFS.scala 673:23]
  wire  _GEN_108 = _T_98 ? 1'h0 : _GEN_102; // @[BFS.scala 695:56 BFS.scala 678:23]
  wire  _GEN_109 = _T_98 ? 1'h0 : _GEN_103; // @[BFS.scala 695:56 BFS.scala 672:28]
  wire [63:0] _GEN_110 = _T_98 ? 64'h0 : _GEN_104; // @[BFS.scala 695:56 BFS.scala 674:25]
  wire [5:0] _GEN_111 = _T_123 ? edge_read_buffer_dout_reg_ptr : _GEN_105; // @[BFS.scala 692:51 BFS.scala 693:23]
  wire  _GEN_112 = _T_123 | _T_98; // @[BFS.scala 692:51 BFS.scala 694:25]
  wire [5:0] _GEN_113 = _T_123 ? 6'h0 : _GEN_107; // @[BFS.scala 692:51 BFS.scala 673:23]
  wire  _GEN_114 = _T_123 ? 1'h0 : _GEN_108; // @[BFS.scala 692:51 BFS.scala 678:23]
  wire  _GEN_115 = _T_123 ? 1'h0 : _GEN_109; // @[BFS.scala 692:51 BFS.scala 672:28]
  wire [63:0] _GEN_116 = _T_123 ? 64'h0 : _GEN_110; // @[BFS.scala 692:51 BFS.scala 674:25]
  wire [5:0] _GEN_117 = _T_120 ? edge_read_buffer_dout_reg_ptr : _GEN_113; // @[BFS.scala 687:55 BFS.scala 688:25]
  wire  _GEN_118 = _T_120 ? _T_116 : _GEN_115; // @[BFS.scala 687:55 BFS.scala 689:30]
  wire [63:0] _GEN_119 = _T_120 ? _num_regfile_io_dataIn_T : _GEN_116; // @[BFS.scala 687:55 BFS.scala 690:27]
  wire [5:0] _GEN_120 = _T_120 ? 6'h0 : _GEN_111; // @[BFS.scala 687:55 BFS.scala 679:21]
  wire  _GEN_121 = _T_120 ? 1'h0 : _GEN_112; // @[BFS.scala 687:55 BFS.scala 680:23]
  wire  _GEN_122 = _T_120 ? 1'h0 : _GEN_114; // @[BFS.scala 687:55 BFS.scala 678:23]
  wire [5:0] _GEN_123 = _T_117 ? free_queue_dout : _GEN_117; // @[BFS.scala 681:46 BFS.scala 682:25]
  wire  _io_read_edge_fifo_empty_T = edge_read_buffer__data_count == 6'h0; // @[util.scala 211:19]
  wire  _credit_dec_T_6 = _T_126 | _T_133; // @[BFS.scala 719:97]
  wire  credit_dec = _credit_dec_T_6 | io_credit_req_valid; // @[BFS.scala 720:82]
  wire  _T_150 = cache_status != 4'h4; // @[BFS.scala 723:18]
  wire  _T_151 = credit_dec & cache_status != 4'h7 & _T_150; // @[BFS.scala 722:63]
  wire [31:0] _credit_T_1 = credit - 32'h1; // @[BFS.scala 724:22]
  wire  _T_156 = ~credit_dec & (_T_122 | _T_123); // @[BFS.scala 725:26]
  wire [31:0] _credit_T_3 = credit + 32'h1; // @[BFS.scala 727:22]
  regFile rid2vid ( // @[BFS.scala 468:23]
    .clock(rid2vid_clock),
    .reset(rid2vid_reset),
    .io_dataIn(rid2vid_io_dataIn),
    .io_dataOut(rid2vid_io_dataOut),
    .io_writeFlag(rid2vid_io_writeFlag),
    .io_rptr(rid2vid_io_rptr),
    .io_wptr(rid2vid_io_wptr)
  );
  regFile_1 num_regfile ( // @[BFS.scala 474:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr)
  );
  meta_fifo edge_read_buffer_ ( // @[BFS.scala 524:32]
    .full(edge_read_buffer__full),
    .din(edge_read_buffer__din),
    .wr_en(edge_read_buffer__wr_en),
    .empty(edge_read_buffer__empty),
    .dout(edge_read_buffer__dout),
    .rd_en(edge_read_buffer__rd_en),
    .data_count(edge_read_buffer__data_count),
    .clk(edge_read_buffer__clk),
    .srst(edge_read_buffer__srst),
    .valid(edge_read_buffer__valid)
  );
  free_queue free_queue ( // @[BFS.scala 574:26]
    .full(free_queue_full),
    .din(free_queue_din),
    .wr_en(free_queue_wr_en),
    .empty(free_queue_empty),
    .dout(free_queue_dout),
    .rd_en(free_queue_rd_en),
    .data_count(free_queue_data_count),
    .clk(free_queue_clk),
    .srst(free_queue_srst),
    .valid(free_queue_valid)
  );
  assign io_in_ready = (~edge_read_buffer__full | status != 2'h0) & io_xbar_out_ready; // @[BFS.scala 555:84]
  assign io_out_valid = _io_out_valid_T_4 | _T_125 | _T_132; // @[BFS.scala 658:89]
  assign io_out_bits_araddr = io_edge_base_addr + _GEN_133; // @[BFS.scala 653:23]
  assign io_out_bits_arid = {1'h1,io_out_bits_arid_lo}; // @[Cat.scala 30:58]
  assign io_out_bits_arlen = arlen[7:0]; // @[BFS.scala 660:21]
  assign io_out_bits_arsize = _io_out_bits_arsize_T ? 3'h2 : _io_out_bits_arsize_T_2; // @[Mux.scala 98:16]
  assign io_xbar_out_valid = io_in_valid & io_in_ready; // @[BFS.scala 515:36]
  assign io_xbar_out_bits_tdata = _T_44 ? _io_xbar_out_bits_tdata_T : io_in_bits_rdata; // @[BFS.scala 517:62 BFS.scala 518:28 BFS.scala 516:26]
  assign io_xbar_out_bits_tkeep = {io_xbar_out_bits_tkeep_hi,io_xbar_out_bits_tkeep_lo}; // @[BFS.scala 521:40]
  assign io_read_edge_fifo_empty = _io_read_edge_fifo_empty_T & _T_105; // @[BFS.scala 717:58]
  assign io_credit = credit[7:0]; // @[BFS.scala 729:13]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 465:21]
  assign rid2vid_clock = clock;
  assign rid2vid_reset = reset;
  assign rid2vid_io_dataIn = io_credit_req_bits_vid; // @[BFS.scala 472:21]
  assign rid2vid_io_writeFlag = io_credit_req_valid; // @[BFS.scala 471:24]
  assign rid2vid_io_rptr = io_in_bits_rid[4:0]; // @[BFS.scala 427:7]
  assign rid2vid_io_wptr = io_credit_req_bits_arid[4:0]; // @[BFS.scala 427:7]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = _T_117 ? _num_regfile_io_dataIn_T : _GEN_119; // @[BFS.scala 681:46 BFS.scala 685:27]
  assign num_regfile_io_writeFlag = _T_117 ? free_queue_valid & io_out_ready & io_out_valid : _GEN_118; // @[BFS.scala 681:46 BFS.scala 684:30]
  assign num_regfile_io_rptr = io_in_bits_rid[4:0]; // @[BFS.scala 427:7]
  assign num_regfile_io_wptr = _GEN_123[4:0];
  assign edge_read_buffer__din = {{1'd0}, _edge_read_buffer_io_din_T}; // @[BFS.scala 535:57]
  assign edge_read_buffer__wr_en = _T_13 & _T; // @[BFS.scala 536:35]
  assign edge_read_buffer__rd_en = cache_status == 4'h9 & init_seq == 6'h0 ? 1'h0 : _GEN_88; // @[BFS.scala 582:60 BFS.scala 534:29]
  assign edge_read_buffer__clk = clock; // @[BFS.scala 527:42]
  assign edge_read_buffer__srst = reset; // @[BFS.scala 528:43]
  assign free_queue_din = _T_117 ? 6'h0 : _GEN_120; // @[BFS.scala 681:46 BFS.scala 679:21]
  assign free_queue_wr_en = _T_117 ? 1'h0 : _GEN_121; // @[BFS.scala 681:46 BFS.scala 680:23]
  assign free_queue_rd_en = _T_117 ? _T_116 : _GEN_122; // @[BFS.scala 681:46 BFS.scala 683:25]
  assign free_queue_clk = clock; // @[BFS.scala 676:36]
  assign free_queue_srst = reset; // @[BFS.scala 677:37]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 445:23]
      status <= 2'h0; // @[BFS.scala 445:23]
    end else if (status == 2'h0 & io_in_valid & io_in_ready) begin // @[BFS.scala 446:63]
      if (io_in_bits_rlast) begin // @[BFS.scala 447:36]
        status <= 2'h0; // @[BFS.scala 448:14]
      end else if (io_in_bits_rid[5]) begin // @[BFS.scala 449:41]
        status <= 2'h2; // @[BFS.scala 450:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 452:14]
      end
    end else if (_T_8 & io_in_valid & io_in_ready & io_in_bits_rlast) begin // @[BFS.scala 455:64]
      status <= 2'h0; // @[BFS.scala 456:12]
    end
    if (reset) begin // @[BFS.scala 458:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 458:35]
    end else if (io_signal) begin // @[BFS.scala 459:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 460:24]
    end else if (_T_17 & _T) begin // @[BFS.scala 462:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 463:24]
    end
    if (reset) begin // @[BFS.scala 475:20]
      num <= 32'h0; // @[BFS.scala 475:20]
    end else if (_T_2 & ~io_in_bits_rlast) begin // @[BFS.scala 477:65]
      if (io_in_bits_rid[5]) begin // @[BFS.scala 478:35]
        if (num_regfile_io_dataOut[63:32] > 32'h4) begin // @[BFS.scala 479:17]
          num <= _num_T_4;
        end else begin
          num <= 32'h0;
        end
      end else if (io_in_bits_rdata[63:32] > 32'h2) begin // @[BFS.scala 481:17]
        num <= _num_T_10;
      end else begin
        num <= 32'h0;
      end
    end else if (_T_6 & io_in_valid & io_in_ready) begin // @[BFS.scala 484:78]
      if (io_in_bits_rlast) begin // @[BFS.scala 485:36]
        num <= 32'h0; // @[BFS.scala 486:11]
      end else begin
        num <= _num_T_13; // @[BFS.scala 488:11]
      end
    end else if (_T_7 & io_in_valid & io_in_ready) begin // @[BFS.scala 490:83]
      num <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 573:29]
      cache_status <= 4'h9; // @[BFS.scala 573:29]
    end else if (cache_status == 4'h9 & init_seq == 6'h0) begin // @[BFS.scala 582:60]
      cache_status <= 4'h6; // @[BFS.scala 583:18]
    end else if (_T_98 & init_seq == 6'h1f) begin // @[BFS.scala 584:77]
      cache_status <= 4'h0; // @[BFS.scala 585:18]
    end else if (cache_status == 4'h0 & edge_read_buffer__valid) begin // @[BFS.scala 586:77]
      cache_status <= {{1'd0}, _GEN_50};
    end else begin
      cache_status <= _GEN_77;
    end
    if (reset) begin // @[BFS.scala 575:25]
      init_seq <= 6'h0; // @[BFS.scala 575:25]
    end else if (cache_status == 4'h6) begin // @[BFS.scala 576:50]
      init_seq <= _init_seq_T_1; // @[BFS.scala 577:14]
    end
    if (reset) begin // @[BFS.scala 579:29]
      expand_index <= 32'h0; // @[BFS.scala 579:29]
    end else if (!(cache_status == 4'h9 & init_seq == 6'h0)) begin // @[BFS.scala 582:60]
      if (!(_T_98 & init_seq == 6'h1f)) begin // @[BFS.scala 584:77]
        if (cache_status == 4'h0 & edge_read_buffer__valid) begin // @[BFS.scala 586:77]
          expand_index <= _GEN_51;
        end else begin
          expand_index <= _GEN_79;
        end
      end
    end
    if (reset) begin // @[BFS.scala 580:29]
      expand_count <= 32'h0; // @[BFS.scala 580:29]
    end else if (!(cache_status == 4'h9 & init_seq == 6'h0)) begin // @[BFS.scala 582:60]
      if (!(_T_98 & init_seq == 6'h1f)) begin // @[BFS.scala 584:77]
        if (cache_status == 4'h0 & edge_read_buffer__valid) begin // @[BFS.scala 586:77]
          expand_count <= _GEN_52;
        end else begin
          expand_count <= _GEN_80;
        end
      end
    end
    if (reset) begin // @[BFS.scala 581:23]
      credit <= 32'h20; // @[BFS.scala 581:23]
    end else if (_T_151) begin // @[BFS.scala 723:42]
      credit <= _credit_T_1; // @[BFS.scala 724:12]
    end else if (_T_156) begin // @[BFS.scala 726:43]
      credit <= _credit_T_3; // @[BFS.scala 727:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  status = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  num = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cache_status = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  init_seq = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  expand_index = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  expand_count = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  credit = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AMBA_Arbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_araddr,
  input  [5:0]  io_in_0_bits_arid,
  input  [7:0]  io_in_0_bits_arlen,
  input  [2:0]  io_in_0_bits_arsize,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_araddr,
  input  [5:0]  io_in_1_bits_arid,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_araddr,
  output [5:0]  io_out_bits_arid,
  output [7:0]  io_out_bits_arlen,
  output [2:0]  io_out_bits_arsize
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  status; // @[util.scala 374:23]
  wire  grant_1 = ~io_in_0_valid; // @[util.scala 363:78]
  reg  grant_reg_0; // @[util.scala 376:26]
  reg  grant_reg_1; // @[util.scala 376:26]
  wire  _T = ~status; // @[util.scala 381:17]
  wire [2:0] _GEN_3 = io_in_0_valid ? io_in_0_bits_arsize : 3'h4; // @[util.scala 382:28 util.scala 384:21 util.scala 379:15]
  wire [7:0] _GEN_4 = io_in_0_valid ? io_in_0_bits_arlen : 8'h3; // @[util.scala 382:28 util.scala 384:21 util.scala 379:15]
  wire [5:0] _GEN_5 = io_in_0_valid ? io_in_0_bits_arid : io_in_1_bits_arid; // @[util.scala 382:28 util.scala 384:21 util.scala 379:15]
  wire [63:0] _GEN_6 = io_in_0_valid ? io_in_0_bits_araddr : io_in_1_bits_araddr; // @[util.scala 382:28 util.scala 384:21 util.scala 379:15]
  wire [2:0] _GEN_10 = grant_reg_0 ? io_in_0_bits_arsize : 3'h4; // @[util.scala 387:26 util.scala 389:21 util.scala 379:15]
  wire [7:0] _GEN_11 = grant_reg_0 ? io_in_0_bits_arlen : 8'h3; // @[util.scala 387:26 util.scala 389:21 util.scala 379:15]
  wire [5:0] _GEN_12 = grant_reg_0 ? io_in_0_bits_arid : io_in_1_bits_arid; // @[util.scala 387:26 util.scala 389:21 util.scala 379:15]
  wire [63:0] _GEN_13 = grant_reg_0 ? io_in_0_bits_araddr : io_in_1_bits_araddr; // @[util.scala 387:26 util.scala 389:21 util.scala 379:15]
  wire [2:0] _GEN_17 = status ? _GEN_10 : 3'h4; // @[util.scala 386:35 util.scala 379:15]
  wire [7:0] _GEN_18 = status ? _GEN_11 : 8'h3; // @[util.scala 386:35 util.scala 379:15]
  wire [5:0] _GEN_19 = status ? _GEN_12 : io_in_1_bits_arid; // @[util.scala 386:35 util.scala 379:15]
  wire [63:0] _GEN_20 = status ? _GEN_13 : io_in_1_bits_araddr; // @[util.scala 386:35 util.scala 379:15]
  wire  _T_8 = grant_1 & io_in_1_valid; // @[util.scala 396:24]
  wire  _GEN_28 = io_out_valid & io_out_ready & status ? 1'h0 : status; // @[util.scala 399:66 util.scala 400:12 util.scala 374:23]
  wire  _GEN_31 = (io_in_0_valid | io_in_1_valid) & _T & ~io_out_ready | _GEN_28; // @[util.scala 394:90 util.scala 398:12]
  assign io_in_0_ready = _T ? io_out_ready : grant_reg_0 & io_out_ready; // @[util.scala 403:20]
  assign io_in_1_ready = _T ? grant_1 & io_out_ready : grant_reg_1 & io_out_ready; // @[util.scala 403:20]
  assign io_out_valid = _T ? ~grant_1 | io_in_1_valid : ~grant_reg_1 | io_in_1_valid; // @[util.scala 405:22]
  assign io_out_bits_araddr = ~status ? _GEN_6 : _GEN_20; // @[util.scala 381:30]
  assign io_out_bits_arid = ~status ? _GEN_5 : _GEN_19; // @[util.scala 381:30]
  assign io_out_bits_arlen = ~status ? _GEN_4 : _GEN_18; // @[util.scala 381:30]
  assign io_out_bits_arsize = ~status ? _GEN_3 : _GEN_17; // @[util.scala 381:30]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 374:23]
      status <= 1'h0; // @[util.scala 374:23]
    end else begin
      status <= _GEN_31;
    end
    if (reset) begin // @[util.scala 376:26]
      grant_reg_0 <= 1'h0; // @[util.scala 376:26]
    end else if ((io_in_0_valid | io_in_1_valid) & _T & ~io_out_ready) begin // @[util.scala 394:90]
      grant_reg_0 <= io_in_0_valid; // @[util.scala 395:15]
    end
    if (reset) begin // @[util.scala 376:26]
      grant_reg_1 <= 1'h0; // @[util.scala 376:26]
    end else if ((io_in_0_valid | io_in_1_valid) & _T & ~io_out_ready) begin // @[util.scala 394:90]
      grant_reg_1 <= _T_8; // @[util.scala 395:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  status = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  grant_reg_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  grant_reg_1 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  output         io_xbar_out_bits_tlast,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  input          io_start,
  input  [31:0]  io_root,
  output         io_issue_sync,
  input  [3:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 770:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 770:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 770:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 770:34]
  wire  edge_cache_clock; // @[BFS.scala 777:26]
  wire  edge_cache_reset; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 777:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 777:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 777:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 777:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 777:26]
  wire  edge_cache_io_xbar_out_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_xbar_out_valid; // @[BFS.scala 777:26]
  wire [127:0] edge_cache_io_xbar_out_bits_tdata; // @[BFS.scala 777:26]
  wire [3:0] edge_cache_io_xbar_out_bits_tkeep; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 777:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 777:26]
  wire [7:0] edge_cache_io_credit; // @[BFS.scala 777:26]
  wire  edge_cache_io_credit_req_valid; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_credit_req_bits_arid; // @[BFS.scala 777:26]
  wire [31:0] edge_cache_io_credit_req_bits_vid; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_traveled_edges; // @[BFS.scala 777:26]
  wire  edge_cache_io_signal; // @[BFS.scala 777:26]
  wire  arbi_clock; // @[BFS.scala 784:20]
  wire  arbi_reset; // @[BFS.scala 784:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 784:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 784:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 784:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 784:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 784:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 784:20]
  wire  arbi_io_out_ready; // @[BFS.scala 784:20]
  wire  arbi_io_out_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 784:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 784:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 784:20]
  wire  vertex_out_fifo_s_axis_aclk; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_aresetn; // @[BFS.scala 813:31]
  wire [127:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 813:31]
  wire [15:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 813:31]
  wire [127:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 813:31]
  wire [15:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 813:31]
  wire [31:0] vertex_out_fifo_axis_rd_data_count; // @[BFS.scala 813:31]
  reg [2:0] upward_status; // @[BFS.scala 766:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 767:30]
  reg [4:0] vertex_read_id; // @[BFS.scala 785:31]
  wire [4:0] _vertex_read_id_T_1 = vertex_read_id + 5'h1; // @[BFS.scala 787:38]
  wire [36:0] _arbi_io_in_1_bits_araddr_T_1 = {vertex_read_buffer_dout[30:0], 6'h0}; // @[BFS.scala 755:59]
  wire [63:0] _GEN_28 = {{27'd0}, _arbi_io_in_1_bits_araddr_T_1}; // @[BFS.scala 755:28]
  wire  _arbi_io_in_1_valid_T_3 = edge_cache_io_credit != 8'h0; // @[BFS.scala 792:26]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 798:104]
  wire  _T_2 = upward_status != 3'h0; // @[BFS.scala 804:88]
  wire  _T_3 = ~io_ddr_r_valid & upward_status != 3'h0; // @[BFS.scala 804:71]
    (*dont_touch = "true" *)reg [30:0] ar_ready_counter; // @[Counter.scala 60:40]
  wire  wrap_wrap = ar_ready_counter == 31'h7ffffffe; // @[Counter.scala 72:24]
  wire [30:0] _wrap_value_T_1 = ar_ready_counter + 31'h1; // @[Counter.scala 76:24]
  wire  _T_6 = io_ddr_r_valid & _T_2; // @[BFS.scala 807:72]
    (*dont_touch = "true" *)reg [30:0] ar_ready_counter_2; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = ar_ready_counter_2 == 31'h7ffffffe; // @[Counter.scala 72:24]
  wire [30:0] _wrap_value_T_3 = ar_ready_counter_2 + 31'h1; // @[Counter.scala 76:24]
  wire [15:0] _io_xbar_out_bits_tkeep_T = vertex_out_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [127:0] _vertex_out_fifo_io_s_axis_tdata_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 128'h80000000 :
    edge_cache_io_xbar_out_bits_tdata; // @[Mux.scala 98:16]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 4'h1 :
    edge_cache_io_xbar_out_bits_tkeep; // @[Mux.scala 98:16]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_2 = io_start ? 4'h1 : _vertex_out_fifo_io_s_axis_tkeep_T_1; // @[Mux.scala 98:16]
  wire  _T_7 = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 831:81]
    (*dont_touch = "true" *)reg [27:0] edge_fifo_ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_5 = edge_fifo_ready_counter + 28'h1; // @[Counter.scala 76:24]
  reg  syncRecv_0; // @[BFS.scala 835:25]
  reg  syncRecv_1; // @[BFS.scala 835:25]
  reg  syncRecv_2; // @[BFS.scala 835:25]
  reg  syncRecv_3; // @[BFS.scala 835:25]
  wire  _GEN_9 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_11 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_13 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_15 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 845:34]
  wire [31:0] _T_15 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_19 = _T_15[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_28 = vertex_out_fifo_axis_rd_data_count == 32'h0; // @[util.scala 320:27]
  wire  _T_29 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_28; // @[BFS.scala 850:71]
  wire [2:0] _GEN_18 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 859:53 BFS.scala 860:19 BFS.scala 766:30]
  wire [2:0] _GEN_19 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3) ? 3'h3 : _GEN_18; // @[BFS.scala 853:71]
  wire  _T_41 = io_xbar_out_valid & ~io_xbar_out_ready; // @[BFS.scala 863:65]
    (*dont_touch = "true" *)reg [27:0] ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_7 = ready_counter + 28'h1; // @[Counter.scala 76:24]
  wire  _T_42 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 866:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 870:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 872:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 770:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 777:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_xbar_out_ready(edge_cache_io_xbar_out_ready),
    .io_xbar_out_valid(edge_cache_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(edge_cache_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(edge_cache_io_xbar_out_bits_tkeep),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_credit(edge_cache_io_credit),
    .io_credit_req_valid(edge_cache_io_credit_req_valid),
    .io_credit_req_bits_arid(edge_cache_io_credit_req_bits_arid),
    .io_credit_req_bits_vid(edge_cache_io_credit_req_bits_vid),
    .io_traveled_edges(edge_cache_io_traveled_edges),
    .io_signal(edge_cache_io_signal)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 784:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 813:31]
    .s_axis_aclk(vertex_out_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_out_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_out_fifo_axis_rd_data_count)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 789:13]
  assign io_ddr_r_ready = edge_cache_io_in_ready; // @[BFS.scala 780:20]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 775:52]
  assign io_xbar_out_valid = vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 817:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_xbar_out_bits_tlast = vertex_out_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_traveled_edges = edge_cache_io_traveled_edges; // @[BFS.scala 781:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 845:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 774:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 773:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 798:88]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 771:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 772:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = io_ddr_r_valid; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rdata = io_ddr_r_bits_rdata; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rid = io_ddr_r_bits_rid; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rlast = io_ddr_r_bits_rlast; // @[BFS.scala 780:20]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 799:17]
  assign edge_cache_io_xbar_out_ready = vertex_out_fifo_s_axis_tready; // @[BFS.scala 829:32]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 779:32]
  assign edge_cache_io_credit_req_valid = arbi_io_in_1_valid & arbi_io_in_1_ready; // @[BFS.scala 800:57]
  assign edge_cache_io_credit_req_bits_arid = arbi_io_in_1_bits_arid; // @[BFS.scala 802:38]
  assign edge_cache_io_credit_req_bits_vid = vertex_read_buffer_dout; // @[BFS.scala 801:37]
  assign edge_cache_io_signal = io_signal; // @[BFS.scala 782:24]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 799:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & _arbi_io_in_1_valid_T_3; // @[BFS.scala 791:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_28; // @[BFS.scala 755:28]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 789:13]
  assign vertex_out_fifo_s_axis_aclk = clock; // @[BFS.scala 815:49]
  assign vertex_out_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 814:40]
  assign vertex_out_fifo_s_axis_tdata = io_start ? {{96'd0}, io_root} : _vertex_out_fifo_io_s_axis_tdata_T_1; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tkeep = {{12'd0}, _vertex_out_fifo_io_s_axis_tkeep_T_2}; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tvalid = edge_cache_io_xbar_out_valid | _vertex_read_buffer_io_rd_en_T_2 | io_start; // @[BFS.scala 819:109]
  assign vertex_out_fifo_s_axis_tlast = 1'h1; // @[BFS.scala 828:35]
  assign vertex_out_fifo_m_axis_tready = io_xbar_out_ready; // @[BFS.scala 818:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 766:30]
      upward_status <= 3'h0; // @[BFS.scala 766:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 846:57]
      upward_status <= 3'h1; // @[BFS.scala 847:19]
    end else if (upward_status == 3'h1 & (_T_19 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3))) begin // @[BFS.scala 848:105]
      upward_status <= 3'h2; // @[BFS.scala 849:19]
    end else if (_T_29 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 851:62]
      upward_status <= 3'h4; // @[BFS.scala 852:19]
    end else begin
      upward_status <= _GEN_19;
    end
    if (reset) begin // @[BFS.scala 767:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 767:30]
    end else if (!(_T_42 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 867:91]
      if (_T_42) begin // @[BFS.scala 869:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 870:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 871:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 872:19]
      end
    end
    if (reset) begin // @[BFS.scala 785:31]
      vertex_read_id <= 5'h0; // @[BFS.scala 785:31]
    end else if (arbi_io_in_1_valid & arbi_io_in_1_ready) begin // @[BFS.scala 786:51]
      vertex_read_id <= _vertex_read_id_T_1; // @[BFS.scala 787:20]
    end
    if (reset) begin // @[Counter.scala 60:40]
      ar_ready_counter <= 31'h0; // @[Counter.scala 60:40]
    end else if (_T_3) begin // @[Counter.scala 118:17]
      if (wrap_wrap) begin // @[Counter.scala 86:20]
        ar_ready_counter <= 31'h0; // @[Counter.scala 86:28]
      end else begin
        ar_ready_counter <= _wrap_value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      ar_ready_counter_2 <= 31'h0; // @[Counter.scala 60:40]
    end else if (_T_6) begin // @[Counter.scala 118:17]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20]
        ar_ready_counter_2 <= 31'h0; // @[Counter.scala 86:28]
      end else begin
        ar_ready_counter_2 <= _wrap_value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      edge_fifo_ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_7) begin // @[Counter.scala 118:17]
      edge_fifo_ready_counter <= _wrap_value_T_5; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_0 <= _GEN_9;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_1 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_2 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_3 <= _GEN_15;
    end
    if (reset) begin // @[Counter.scala 60:40]
      ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_41) begin // @[Counter.scala 118:17]
      ready_counter <= _wrap_value_T_7; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  vertex_read_id = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  ar_ready_counter = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  ar_ready_counter_2 = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  edge_fifo_ready_counter = _RAND_5[27:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  syncRecv_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_1(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  output         io_xbar_out_bits_tlast,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [3:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 770:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 770:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 770:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 770:34]
  wire  edge_cache_clock; // @[BFS.scala 777:26]
  wire  edge_cache_reset; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 777:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 777:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 777:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 777:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 777:26]
  wire  edge_cache_io_xbar_out_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_xbar_out_valid; // @[BFS.scala 777:26]
  wire [127:0] edge_cache_io_xbar_out_bits_tdata; // @[BFS.scala 777:26]
  wire [3:0] edge_cache_io_xbar_out_bits_tkeep; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 777:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 777:26]
  wire [7:0] edge_cache_io_credit; // @[BFS.scala 777:26]
  wire  edge_cache_io_credit_req_valid; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_credit_req_bits_arid; // @[BFS.scala 777:26]
  wire [31:0] edge_cache_io_credit_req_bits_vid; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_traveled_edges; // @[BFS.scala 777:26]
  wire  edge_cache_io_signal; // @[BFS.scala 777:26]
  wire  arbi_clock; // @[BFS.scala 784:20]
  wire  arbi_reset; // @[BFS.scala 784:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 784:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 784:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 784:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 784:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 784:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 784:20]
  wire  arbi_io_out_ready; // @[BFS.scala 784:20]
  wire  arbi_io_out_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 784:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 784:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 784:20]
  wire  vertex_out_fifo_s_axis_aclk; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_aresetn; // @[BFS.scala 813:31]
  wire [127:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 813:31]
  wire [15:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 813:31]
  wire [127:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 813:31]
  wire [15:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 813:31]
  wire [31:0] vertex_out_fifo_axis_rd_data_count; // @[BFS.scala 813:31]
  reg [2:0] upward_status; // @[BFS.scala 766:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 767:30]
  reg [4:0] vertex_read_id; // @[BFS.scala 785:31]
  wire [4:0] _vertex_read_id_T_1 = vertex_read_id + 5'h1; // @[BFS.scala 787:38]
  wire [36:0] _arbi_io_in_1_bits_araddr_T_1 = {vertex_read_buffer_dout[30:0], 6'h0}; // @[BFS.scala 755:59]
  wire [63:0] _GEN_28 = {{27'd0}, _arbi_io_in_1_bits_araddr_T_1}; // @[BFS.scala 755:28]
  wire  _arbi_io_in_1_valid_T_3 = edge_cache_io_credit != 8'h0; // @[BFS.scala 792:26]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 798:104]
  wire  _T_2 = upward_status != 3'h0; // @[BFS.scala 804:88]
  wire  _T_3 = ~io_ddr_r_valid & upward_status != 3'h0; // @[BFS.scala 804:71]
    (*dont_touch = "true" *)reg [30:0] ar_ready_counter; // @[Counter.scala 60:40]
  wire  wrap_wrap = ar_ready_counter == 31'h7ffffffe; // @[Counter.scala 72:24]
  wire [30:0] _wrap_value_T_1 = ar_ready_counter + 31'h1; // @[Counter.scala 76:24]
  wire  _T_6 = io_ddr_r_valid & _T_2; // @[BFS.scala 807:72]
    (*dont_touch = "true" *)reg [30:0] ar_ready_counter_2; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = ar_ready_counter_2 == 31'h7ffffffe; // @[Counter.scala 72:24]
  wire [30:0] _wrap_value_T_3 = ar_ready_counter_2 + 31'h1; // @[Counter.scala 76:24]
  wire [15:0] _io_xbar_out_bits_tkeep_T = vertex_out_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 4'h1 :
    edge_cache_io_xbar_out_bits_tkeep; // @[Mux.scala 98:16]
  wire  _T_7 = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 831:81]
    (*dont_touch = "true" *)reg [27:0] edge_fifo_ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_5 = edge_fifo_ready_counter + 28'h1; // @[Counter.scala 76:24]
  reg  syncRecv_0; // @[BFS.scala 835:25]
  reg  syncRecv_1; // @[BFS.scala 835:25]
  reg  syncRecv_2; // @[BFS.scala 835:25]
  reg  syncRecv_3; // @[BFS.scala 835:25]
  wire  _GEN_9 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_11 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_13 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_15 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 845:34]
  wire [31:0] _T_15 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_19 = _T_15[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_28 = vertex_out_fifo_axis_rd_data_count == 32'h0; // @[util.scala 320:27]
  wire  _T_29 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_28; // @[BFS.scala 850:71]
  wire [2:0] _GEN_18 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 859:53 BFS.scala 860:19 BFS.scala 766:30]
  wire [2:0] _GEN_19 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3) ? 3'h0 : _GEN_18; // @[BFS.scala 853:71]
  wire  _T_41 = io_xbar_out_valid & ~io_xbar_out_ready; // @[BFS.scala 863:65]
    (*dont_touch = "true" *)reg [27:0] ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_7 = ready_counter + 28'h1; // @[Counter.scala 76:24]
  wire  _T_42 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 866:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 870:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 872:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 770:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 777:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_xbar_out_ready(edge_cache_io_xbar_out_ready),
    .io_xbar_out_valid(edge_cache_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(edge_cache_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(edge_cache_io_xbar_out_bits_tkeep),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_credit(edge_cache_io_credit),
    .io_credit_req_valid(edge_cache_io_credit_req_valid),
    .io_credit_req_bits_arid(edge_cache_io_credit_req_bits_arid),
    .io_credit_req_bits_vid(edge_cache_io_credit_req_bits_vid),
    .io_traveled_edges(edge_cache_io_traveled_edges),
    .io_signal(edge_cache_io_signal)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 784:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 813:31]
    .s_axis_aclk(vertex_out_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_out_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_out_fifo_axis_rd_data_count)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 789:13]
  assign io_ddr_r_ready = edge_cache_io_in_ready; // @[BFS.scala 780:20]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 775:52]
  assign io_xbar_out_valid = vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 817:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_xbar_out_bits_tlast = vertex_out_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_traveled_edges = edge_cache_io_traveled_edges; // @[BFS.scala 781:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 845:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 774:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 773:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 798:88]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 771:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 772:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = io_ddr_r_valid; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rdata = io_ddr_r_bits_rdata; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rid = io_ddr_r_bits_rid; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rlast = io_ddr_r_bits_rlast; // @[BFS.scala 780:20]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 799:17]
  assign edge_cache_io_xbar_out_ready = vertex_out_fifo_s_axis_tready; // @[BFS.scala 829:32]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 779:32]
  assign edge_cache_io_credit_req_valid = arbi_io_in_1_valid & arbi_io_in_1_ready; // @[BFS.scala 800:57]
  assign edge_cache_io_credit_req_bits_arid = arbi_io_in_1_bits_arid; // @[BFS.scala 802:38]
  assign edge_cache_io_credit_req_bits_vid = vertex_read_buffer_dout; // @[BFS.scala 801:37]
  assign edge_cache_io_signal = io_signal; // @[BFS.scala 782:24]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 799:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & _arbi_io_in_1_valid_T_3; // @[BFS.scala 791:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_28; // @[BFS.scala 755:28]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 789:13]
  assign vertex_out_fifo_s_axis_aclk = clock; // @[BFS.scala 815:49]
  assign vertex_out_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 814:40]
  assign vertex_out_fifo_s_axis_tdata = _vertex_read_buffer_io_rd_en_T_2 ? 128'h80000000 :
    edge_cache_io_xbar_out_bits_tdata; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tkeep = {{12'd0}, _vertex_out_fifo_io_s_axis_tkeep_T_1}; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tvalid = edge_cache_io_xbar_out_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 819:68]
  assign vertex_out_fifo_s_axis_tlast = 1'h1; // @[BFS.scala 828:35]
  assign vertex_out_fifo_m_axis_tready = io_xbar_out_ready; // @[BFS.scala 818:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 766:30]
      upward_status <= 3'h0; // @[BFS.scala 766:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 846:57]
      upward_status <= 3'h1; // @[BFS.scala 847:19]
    end else if (upward_status == 3'h1 & (_T_19 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3))) begin // @[BFS.scala 848:105]
      upward_status <= 3'h2; // @[BFS.scala 849:19]
    end else if (_T_29 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 851:62]
      upward_status <= 3'h4; // @[BFS.scala 852:19]
    end else begin
      upward_status <= _GEN_19;
    end
    if (reset) begin // @[BFS.scala 767:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 767:30]
    end else if (!(_T_42 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 867:91]
      if (_T_42) begin // @[BFS.scala 869:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 870:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 871:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 872:19]
      end
    end
    if (reset) begin // @[BFS.scala 785:31]
      vertex_read_id <= 5'h0; // @[BFS.scala 785:31]
    end else if (arbi_io_in_1_valid & arbi_io_in_1_ready) begin // @[BFS.scala 786:51]
      vertex_read_id <= _vertex_read_id_T_1; // @[BFS.scala 787:20]
    end
    if (reset) begin // @[Counter.scala 60:40]
      ar_ready_counter <= 31'h0; // @[Counter.scala 60:40]
    end else if (_T_3) begin // @[Counter.scala 118:17]
      if (wrap_wrap) begin // @[Counter.scala 86:20]
        ar_ready_counter <= 31'h0; // @[Counter.scala 86:28]
      end else begin
        ar_ready_counter <= _wrap_value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      ar_ready_counter_2 <= 31'h0; // @[Counter.scala 60:40]
    end else if (_T_6) begin // @[Counter.scala 118:17]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20]
        ar_ready_counter_2 <= 31'h0; // @[Counter.scala 86:28]
      end else begin
        ar_ready_counter_2 <= _wrap_value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      edge_fifo_ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_7) begin // @[Counter.scala 118:17]
      edge_fifo_ready_counter <= _wrap_value_T_5; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_0 <= _GEN_9;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_1 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_2 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_3 <= _GEN_15;
    end
    if (reset) begin // @[Counter.scala 60:40]
      ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_41) begin // @[Counter.scala 118:17]
      ready_counter <= _wrap_value_T_7; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  vertex_read_id = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  ar_ready_counter = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  ar_ready_counter_2 = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  edge_fifo_ready_counter = _RAND_5[27:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  syncRecv_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_2(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  output         io_xbar_out_bits_tlast,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [3:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 770:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 770:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 770:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 770:34]
  wire  edge_cache_clock; // @[BFS.scala 777:26]
  wire  edge_cache_reset; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 777:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 777:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 777:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 777:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 777:26]
  wire  edge_cache_io_xbar_out_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_xbar_out_valid; // @[BFS.scala 777:26]
  wire [127:0] edge_cache_io_xbar_out_bits_tdata; // @[BFS.scala 777:26]
  wire [3:0] edge_cache_io_xbar_out_bits_tkeep; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 777:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 777:26]
  wire [7:0] edge_cache_io_credit; // @[BFS.scala 777:26]
  wire  edge_cache_io_credit_req_valid; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_credit_req_bits_arid; // @[BFS.scala 777:26]
  wire [31:0] edge_cache_io_credit_req_bits_vid; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_traveled_edges; // @[BFS.scala 777:26]
  wire  edge_cache_io_signal; // @[BFS.scala 777:26]
  wire  arbi_clock; // @[BFS.scala 784:20]
  wire  arbi_reset; // @[BFS.scala 784:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 784:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 784:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 784:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 784:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 784:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 784:20]
  wire  arbi_io_out_ready; // @[BFS.scala 784:20]
  wire  arbi_io_out_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 784:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 784:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 784:20]
  wire  vertex_out_fifo_s_axis_aclk; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_aresetn; // @[BFS.scala 813:31]
  wire [127:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 813:31]
  wire [15:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 813:31]
  wire [127:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 813:31]
  wire [15:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 813:31]
  wire [31:0] vertex_out_fifo_axis_rd_data_count; // @[BFS.scala 813:31]
  reg [2:0] upward_status; // @[BFS.scala 766:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 767:30]
  reg [4:0] vertex_read_id; // @[BFS.scala 785:31]
  wire [4:0] _vertex_read_id_T_1 = vertex_read_id + 5'h1; // @[BFS.scala 787:38]
  wire [36:0] _arbi_io_in_1_bits_araddr_T_1 = {vertex_read_buffer_dout[30:0], 6'h0}; // @[BFS.scala 755:59]
  wire [63:0] _GEN_28 = {{27'd0}, _arbi_io_in_1_bits_araddr_T_1}; // @[BFS.scala 755:28]
  wire  _arbi_io_in_1_valid_T_3 = edge_cache_io_credit != 8'h0; // @[BFS.scala 792:26]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 798:104]
  wire  _T_2 = upward_status != 3'h0; // @[BFS.scala 804:88]
  wire  _T_3 = ~io_ddr_r_valid & upward_status != 3'h0; // @[BFS.scala 804:71]
    (*dont_touch = "true" *)reg [30:0] ar_ready_counter; // @[Counter.scala 60:40]
  wire  wrap_wrap = ar_ready_counter == 31'h7ffffffe; // @[Counter.scala 72:24]
  wire [30:0] _wrap_value_T_1 = ar_ready_counter + 31'h1; // @[Counter.scala 76:24]
  wire  _T_6 = io_ddr_r_valid & _T_2; // @[BFS.scala 807:72]
    (*dont_touch = "true" *)reg [30:0] ar_ready_counter_2; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = ar_ready_counter_2 == 31'h7ffffffe; // @[Counter.scala 72:24]
  wire [30:0] _wrap_value_T_3 = ar_ready_counter_2 + 31'h1; // @[Counter.scala 76:24]
  wire [15:0] _io_xbar_out_bits_tkeep_T = vertex_out_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 4'h1 :
    edge_cache_io_xbar_out_bits_tkeep; // @[Mux.scala 98:16]
  wire  _T_7 = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 831:81]
    (*dont_touch = "true" *)reg [27:0] edge_fifo_ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_5 = edge_fifo_ready_counter + 28'h1; // @[Counter.scala 76:24]
  reg  syncRecv_0; // @[BFS.scala 835:25]
  reg  syncRecv_1; // @[BFS.scala 835:25]
  reg  syncRecv_2; // @[BFS.scala 835:25]
  reg  syncRecv_3; // @[BFS.scala 835:25]
  wire  _GEN_9 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_11 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_13 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_15 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 845:34]
  wire [31:0] _T_15 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_19 = _T_15[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_28 = vertex_out_fifo_axis_rd_data_count == 32'h0; // @[util.scala 320:27]
  wire  _T_29 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_28; // @[BFS.scala 850:71]
  wire [2:0] _GEN_18 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 859:53 BFS.scala 860:19 BFS.scala 766:30]
  wire [2:0] _GEN_19 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3) ? 3'h0 : _GEN_18; // @[BFS.scala 853:71]
  wire  _T_41 = io_xbar_out_valid & ~io_xbar_out_ready; // @[BFS.scala 863:65]
    (*dont_touch = "true" *)reg [27:0] ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_7 = ready_counter + 28'h1; // @[Counter.scala 76:24]
  wire  _T_42 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 866:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 870:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 872:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 770:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 777:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_xbar_out_ready(edge_cache_io_xbar_out_ready),
    .io_xbar_out_valid(edge_cache_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(edge_cache_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(edge_cache_io_xbar_out_bits_tkeep),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_credit(edge_cache_io_credit),
    .io_credit_req_valid(edge_cache_io_credit_req_valid),
    .io_credit_req_bits_arid(edge_cache_io_credit_req_bits_arid),
    .io_credit_req_bits_vid(edge_cache_io_credit_req_bits_vid),
    .io_traveled_edges(edge_cache_io_traveled_edges),
    .io_signal(edge_cache_io_signal)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 784:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 813:31]
    .s_axis_aclk(vertex_out_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_out_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_out_fifo_axis_rd_data_count)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 789:13]
  assign io_ddr_r_ready = edge_cache_io_in_ready; // @[BFS.scala 780:20]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 775:52]
  assign io_xbar_out_valid = vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 817:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_xbar_out_bits_tlast = vertex_out_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_traveled_edges = edge_cache_io_traveled_edges; // @[BFS.scala 781:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 845:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 774:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 773:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 798:88]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 771:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 772:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = io_ddr_r_valid; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rdata = io_ddr_r_bits_rdata; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rid = io_ddr_r_bits_rid; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rlast = io_ddr_r_bits_rlast; // @[BFS.scala 780:20]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 799:17]
  assign edge_cache_io_xbar_out_ready = vertex_out_fifo_s_axis_tready; // @[BFS.scala 829:32]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 779:32]
  assign edge_cache_io_credit_req_valid = arbi_io_in_1_valid & arbi_io_in_1_ready; // @[BFS.scala 800:57]
  assign edge_cache_io_credit_req_bits_arid = arbi_io_in_1_bits_arid; // @[BFS.scala 802:38]
  assign edge_cache_io_credit_req_bits_vid = vertex_read_buffer_dout; // @[BFS.scala 801:37]
  assign edge_cache_io_signal = io_signal; // @[BFS.scala 782:24]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 799:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & _arbi_io_in_1_valid_T_3; // @[BFS.scala 791:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_28; // @[BFS.scala 755:28]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 789:13]
  assign vertex_out_fifo_s_axis_aclk = clock; // @[BFS.scala 815:49]
  assign vertex_out_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 814:40]
  assign vertex_out_fifo_s_axis_tdata = _vertex_read_buffer_io_rd_en_T_2 ? 128'h80000000 :
    edge_cache_io_xbar_out_bits_tdata; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tkeep = {{12'd0}, _vertex_out_fifo_io_s_axis_tkeep_T_1}; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tvalid = edge_cache_io_xbar_out_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 819:68]
  assign vertex_out_fifo_s_axis_tlast = 1'h1; // @[BFS.scala 828:35]
  assign vertex_out_fifo_m_axis_tready = io_xbar_out_ready; // @[BFS.scala 818:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 766:30]
      upward_status <= 3'h0; // @[BFS.scala 766:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 846:57]
      upward_status <= 3'h1; // @[BFS.scala 847:19]
    end else if (upward_status == 3'h1 & (_T_19 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3))) begin // @[BFS.scala 848:105]
      upward_status <= 3'h2; // @[BFS.scala 849:19]
    end else if (_T_29 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 851:62]
      upward_status <= 3'h4; // @[BFS.scala 852:19]
    end else begin
      upward_status <= _GEN_19;
    end
    if (reset) begin // @[BFS.scala 767:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 767:30]
    end else if (!(_T_42 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 867:91]
      if (_T_42) begin // @[BFS.scala 869:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 870:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 871:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 872:19]
      end
    end
    if (reset) begin // @[BFS.scala 785:31]
      vertex_read_id <= 5'h0; // @[BFS.scala 785:31]
    end else if (arbi_io_in_1_valid & arbi_io_in_1_ready) begin // @[BFS.scala 786:51]
      vertex_read_id <= _vertex_read_id_T_1; // @[BFS.scala 787:20]
    end
    if (reset) begin // @[Counter.scala 60:40]
      ar_ready_counter <= 31'h0; // @[Counter.scala 60:40]
    end else if (_T_3) begin // @[Counter.scala 118:17]
      if (wrap_wrap) begin // @[Counter.scala 86:20]
        ar_ready_counter <= 31'h0; // @[Counter.scala 86:28]
      end else begin
        ar_ready_counter <= _wrap_value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      ar_ready_counter_2 <= 31'h0; // @[Counter.scala 60:40]
    end else if (_T_6) begin // @[Counter.scala 118:17]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20]
        ar_ready_counter_2 <= 31'h0; // @[Counter.scala 86:28]
      end else begin
        ar_ready_counter_2 <= _wrap_value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      edge_fifo_ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_7) begin // @[Counter.scala 118:17]
      edge_fifo_ready_counter <= _wrap_value_T_5; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_0 <= _GEN_9;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_1 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_2 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_3 <= _GEN_15;
    end
    if (reset) begin // @[Counter.scala 60:40]
      ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_41) begin // @[Counter.scala 118:17]
      ready_counter <= _wrap_value_T_7; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  vertex_read_id = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  ar_ready_counter = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  ar_ready_counter_2 = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  edge_fifo_ready_counter = _RAND_5[27:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  syncRecv_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_3(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  output         io_xbar_out_bits_tlast,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [3:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 770:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 770:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 770:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 770:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 770:34]
  wire  edge_cache_clock; // @[BFS.scala 777:26]
  wire  edge_cache_reset; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 777:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 777:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 777:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 777:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 777:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 777:26]
  wire  edge_cache_io_xbar_out_ready; // @[BFS.scala 777:26]
  wire  edge_cache_io_xbar_out_valid; // @[BFS.scala 777:26]
  wire [127:0] edge_cache_io_xbar_out_bits_tdata; // @[BFS.scala 777:26]
  wire [3:0] edge_cache_io_xbar_out_bits_tkeep; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 777:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 777:26]
  wire [7:0] edge_cache_io_credit; // @[BFS.scala 777:26]
  wire  edge_cache_io_credit_req_valid; // @[BFS.scala 777:26]
  wire [5:0] edge_cache_io_credit_req_bits_arid; // @[BFS.scala 777:26]
  wire [31:0] edge_cache_io_credit_req_bits_vid; // @[BFS.scala 777:26]
  wire [63:0] edge_cache_io_traveled_edges; // @[BFS.scala 777:26]
  wire  edge_cache_io_signal; // @[BFS.scala 777:26]
  wire  arbi_clock; // @[BFS.scala 784:20]
  wire  arbi_reset; // @[BFS.scala 784:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 784:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 784:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 784:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 784:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 784:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 784:20]
  wire  arbi_io_out_ready; // @[BFS.scala 784:20]
  wire  arbi_io_out_valid; // @[BFS.scala 784:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 784:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 784:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 784:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 784:20]
  wire  vertex_out_fifo_s_axis_aclk; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_aresetn; // @[BFS.scala 813:31]
  wire [127:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 813:31]
  wire [15:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 813:31]
  wire [127:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 813:31]
  wire [15:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 813:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 813:31]
  wire [31:0] vertex_out_fifo_axis_rd_data_count; // @[BFS.scala 813:31]
  reg [2:0] upward_status; // @[BFS.scala 766:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 767:30]
  reg [4:0] vertex_read_id; // @[BFS.scala 785:31]
  wire [4:0] _vertex_read_id_T_1 = vertex_read_id + 5'h1; // @[BFS.scala 787:38]
  wire [36:0] _arbi_io_in_1_bits_araddr_T_1 = {vertex_read_buffer_dout[30:0], 6'h0}; // @[BFS.scala 755:59]
  wire [63:0] _GEN_28 = {{27'd0}, _arbi_io_in_1_bits_araddr_T_1}; // @[BFS.scala 755:28]
  wire  _arbi_io_in_1_valid_T_3 = edge_cache_io_credit != 8'h0; // @[BFS.scala 792:26]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 798:104]
  wire  _T_2 = upward_status != 3'h0; // @[BFS.scala 804:88]
  wire  _T_3 = ~io_ddr_r_valid & upward_status != 3'h0; // @[BFS.scala 804:71]
    (*dont_touch = "true" *)reg [30:0] ar_ready_counter; // @[Counter.scala 60:40]
  wire  wrap_wrap = ar_ready_counter == 31'h7ffffffe; // @[Counter.scala 72:24]
  wire [30:0] _wrap_value_T_1 = ar_ready_counter + 31'h1; // @[Counter.scala 76:24]
  wire  _T_6 = io_ddr_r_valid & _T_2; // @[BFS.scala 807:72]
    (*dont_touch = "true" *)reg [30:0] ar_ready_counter_2; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = ar_ready_counter_2 == 31'h7ffffffe; // @[Counter.scala 72:24]
  wire [30:0] _wrap_value_T_3 = ar_ready_counter_2 + 31'h1; // @[Counter.scala 76:24]
  wire [15:0] _io_xbar_out_bits_tkeep_T = vertex_out_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 4'h1 :
    edge_cache_io_xbar_out_bits_tkeep; // @[Mux.scala 98:16]
  wire  _T_7 = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 831:81]
    (*dont_touch = "true" *)reg [27:0] edge_fifo_ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_5 = edge_fifo_ready_counter + 28'h1; // @[Counter.scala 76:24]
  reg  syncRecv_0; // @[BFS.scala 835:25]
  reg  syncRecv_1; // @[BFS.scala 835:25]
  reg  syncRecv_2; // @[BFS.scala 835:25]
  reg  syncRecv_3; // @[BFS.scala 835:25]
  wire  _GEN_9 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_11 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_13 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _GEN_15 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 840:34 BFS.scala 841:11 BFS.scala 835:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 845:34]
  wire [31:0] _T_15 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_19 = _T_15[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_28 = vertex_out_fifo_axis_rd_data_count == 32'h0; // @[util.scala 320:27]
  wire  _T_29 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_28; // @[BFS.scala 850:71]
  wire [2:0] _GEN_18 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 859:53 BFS.scala 860:19 BFS.scala 766:30]
  wire [2:0] _GEN_19 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3) ? 3'h0 : _GEN_18; // @[BFS.scala 853:71]
  wire  _T_41 = io_xbar_out_valid & ~io_xbar_out_ready; // @[BFS.scala 863:65]
    (*dont_touch = "true" *)reg [27:0] ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_7 = ready_counter + 28'h1; // @[Counter.scala 76:24]
  wire  _T_42 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 866:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 870:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 872:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 770:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 777:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_xbar_out_ready(edge_cache_io_xbar_out_ready),
    .io_xbar_out_valid(edge_cache_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(edge_cache_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(edge_cache_io_xbar_out_bits_tkeep),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_credit(edge_cache_io_credit),
    .io_credit_req_valid(edge_cache_io_credit_req_valid),
    .io_credit_req_bits_arid(edge_cache_io_credit_req_bits_arid),
    .io_credit_req_bits_vid(edge_cache_io_credit_req_bits_vid),
    .io_traveled_edges(edge_cache_io_traveled_edges),
    .io_signal(edge_cache_io_signal)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 784:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 813:31]
    .s_axis_aclk(vertex_out_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_out_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_out_fifo_axis_rd_data_count)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 789:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 789:13]
  assign io_ddr_r_ready = edge_cache_io_in_ready; // @[BFS.scala 780:20]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 775:52]
  assign io_xbar_out_valid = vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 817:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_xbar_out_bits_tlast = vertex_out_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_traveled_edges = edge_cache_io_traveled_edges; // @[BFS.scala 781:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 845:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 774:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 773:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 798:88]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 771:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 772:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = io_ddr_r_valid; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rdata = io_ddr_r_bits_rdata; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rid = io_ddr_r_bits_rid; // @[BFS.scala 780:20]
  assign edge_cache_io_in_bits_rlast = io_ddr_r_bits_rlast; // @[BFS.scala 780:20]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 799:17]
  assign edge_cache_io_xbar_out_ready = vertex_out_fifo_s_axis_tready; // @[BFS.scala 829:32]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 779:32]
  assign edge_cache_io_credit_req_valid = arbi_io_in_1_valid & arbi_io_in_1_ready; // @[BFS.scala 800:57]
  assign edge_cache_io_credit_req_bits_arid = arbi_io_in_1_bits_arid; // @[BFS.scala 802:38]
  assign edge_cache_io_credit_req_bits_vid = vertex_read_buffer_dout; // @[BFS.scala 801:37]
  assign edge_cache_io_signal = io_signal; // @[BFS.scala 782:24]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 799:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 799:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & _arbi_io_in_1_valid_T_3; // @[BFS.scala 791:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_28; // @[BFS.scala 755:28]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 789:13]
  assign vertex_out_fifo_s_axis_aclk = clock; // @[BFS.scala 815:49]
  assign vertex_out_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 814:40]
  assign vertex_out_fifo_s_axis_tdata = _vertex_read_buffer_io_rd_en_T_2 ? 128'h80000000 :
    edge_cache_io_xbar_out_bits_tdata; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tkeep = {{12'd0}, _vertex_out_fifo_io_s_axis_tkeep_T_1}; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tvalid = edge_cache_io_xbar_out_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 819:68]
  assign vertex_out_fifo_s_axis_tlast = 1'h1; // @[BFS.scala 828:35]
  assign vertex_out_fifo_m_axis_tready = io_xbar_out_ready; // @[BFS.scala 818:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 766:30]
      upward_status <= 3'h0; // @[BFS.scala 766:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 846:57]
      upward_status <= 3'h1; // @[BFS.scala 847:19]
    end else if (upward_status == 3'h1 & (_T_19 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3))) begin // @[BFS.scala 848:105]
      upward_status <= 3'h2; // @[BFS.scala 849:19]
    end else if (_T_29 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 851:62]
      upward_status <= 3'h4; // @[BFS.scala 852:19]
    end else begin
      upward_status <= _GEN_19;
    end
    if (reset) begin // @[BFS.scala 767:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 767:30]
    end else if (!(_T_42 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 867:91]
      if (_T_42) begin // @[BFS.scala 869:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 870:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 871:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 872:19]
      end
    end
    if (reset) begin // @[BFS.scala 785:31]
      vertex_read_id <= 5'h0; // @[BFS.scala 785:31]
    end else if (arbi_io_in_1_valid & arbi_io_in_1_ready) begin // @[BFS.scala 786:51]
      vertex_read_id <= _vertex_read_id_T_1; // @[BFS.scala 787:20]
    end
    if (reset) begin // @[Counter.scala 60:40]
      ar_ready_counter <= 31'h0; // @[Counter.scala 60:40]
    end else if (_T_3) begin // @[Counter.scala 118:17]
      if (wrap_wrap) begin // @[Counter.scala 86:20]
        ar_ready_counter <= 31'h0; // @[Counter.scala 86:28]
      end else begin
        ar_ready_counter <= _wrap_value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      ar_ready_counter_2 <= 31'h0; // @[Counter.scala 60:40]
    end else if (_T_6) begin // @[Counter.scala 118:17]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20]
        ar_ready_counter_2 <= 31'h0; // @[Counter.scala 86:28]
      end else begin
        ar_ready_counter_2 <= _wrap_value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      edge_fifo_ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_7) begin // @[Counter.scala 118:17]
      edge_fifo_ready_counter <= _wrap_value_T_5; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_0 <= _GEN_9;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_1 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_2 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 835:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 835:25]
    end else if (io_signal) begin // @[BFS.scala 838:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 839:11]
    end else begin
      syncRecv_3 <= _GEN_15;
    end
    if (reset) begin // @[Counter.scala 60:40]
      ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_41) begin // @[Counter.scala 118:17]
      ready_counter <= _wrap_value_T_7; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  vertex_read_id = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  ar_ready_counter = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  ar_ready_counter_2 = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  edge_fifo_ready_counter = _RAND_5[27:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  syncRecv_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fat_vertex_cache(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [511:0] io_ddr_out_bits_tdata,
  output [15:0]  io_ddr_out_bits_tkeep,
  output         io_ddr_out_bits_tlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  filter_0_aclk; // @[BFS.scala 882:34]
  wire  filter_0_aresetn; // @[BFS.scala 882:34]
  wire [511:0] filter_0_s_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_0_s_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_0_s_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_0_s_axis_tready; // @[BFS.scala 882:34]
  wire  filter_0_s_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_0_s_axis_tuser; // @[BFS.scala 882:34]
  wire [511:0] filter_0_m_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_0_m_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_0_m_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_0_m_axis_tready; // @[BFS.scala 882:34]
  wire  filter_0_m_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_0_m_axis_tuser; // @[BFS.scala 882:34]
  wire  filter_1_aclk; // @[BFS.scala 882:34]
  wire  filter_1_aresetn; // @[BFS.scala 882:34]
  wire [511:0] filter_1_s_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_1_s_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_1_s_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_1_s_axis_tready; // @[BFS.scala 882:34]
  wire  filter_1_s_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_1_s_axis_tuser; // @[BFS.scala 882:34]
  wire [511:0] filter_1_m_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_1_m_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_1_m_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_1_m_axis_tready; // @[BFS.scala 882:34]
  wire  filter_1_m_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_1_m_axis_tuser; // @[BFS.scala 882:34]
  wire  filter_2_aclk; // @[BFS.scala 882:34]
  wire  filter_2_aresetn; // @[BFS.scala 882:34]
  wire [511:0] filter_2_s_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_2_s_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_2_s_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_2_s_axis_tready; // @[BFS.scala 882:34]
  wire  filter_2_s_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_2_s_axis_tuser; // @[BFS.scala 882:34]
  wire [511:0] filter_2_m_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_2_m_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_2_m_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_2_m_axis_tready; // @[BFS.scala 882:34]
  wire  filter_2_m_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_2_m_axis_tuser; // @[BFS.scala 882:34]
  wire  filter_3_aclk; // @[BFS.scala 882:34]
  wire  filter_3_aresetn; // @[BFS.scala 882:34]
  wire [511:0] filter_3_s_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_3_s_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_3_s_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_3_s_axis_tready; // @[BFS.scala 882:34]
  wire  filter_3_s_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_3_s_axis_tuser; // @[BFS.scala 882:34]
  wire [511:0] filter_3_m_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_3_m_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_3_m_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_3_m_axis_tready; // @[BFS.scala 882:34]
  wire  filter_3_m_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_3_m_axis_tuser; // @[BFS.scala 882:34]
  wire  filter_4_aclk; // @[BFS.scala 882:34]
  wire  filter_4_aresetn; // @[BFS.scala 882:34]
  wire [511:0] filter_4_s_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_4_s_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_4_s_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_4_s_axis_tready; // @[BFS.scala 882:34]
  wire  filter_4_s_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_4_s_axis_tuser; // @[BFS.scala 882:34]
  wire [511:0] filter_4_m_axis_tdata; // @[BFS.scala 882:34]
  wire [63:0] filter_4_m_axis_tkeep; // @[BFS.scala 882:34]
  wire  filter_4_m_axis_tvalid; // @[BFS.scala 882:34]
  wire  filter_4_m_axis_tready; // @[BFS.scala 882:34]
  wire  filter_4_m_axis_tlast; // @[BFS.scala 882:34]
  wire [3:0] filter_4_m_axis_tuser; // @[BFS.scala 882:34]
  reg  fat_vertex_entry_0_valid; // @[BFS.scala 884:46]
  reg [63:0] fat_vertex_entry_0_bits; // @[BFS.scala 884:46]
  reg  fat_vertex_entry_1_valid; // @[BFS.scala 884:46]
  reg [63:0] fat_vertex_entry_1_bits; // @[BFS.scala 884:46]
  reg  fat_vertex_entry_2_valid; // @[BFS.scala 884:46]
  reg [63:0] fat_vertex_entry_2_bits; // @[BFS.scala 884:46]
  reg  fat_vertex_entry_3_valid; // @[BFS.scala 884:46]
  reg [63:0] fat_vertex_entry_3_bits; // @[BFS.scala 884:46]
  wire [1:0] filter_0_io_s_axis_tuser_lo = {io_xbar_in_bits_tkeep[6:4] == 3'h4,io_xbar_in_bits_tkeep[2:0] == 3'h4}; // @[BFS.scala 886:106]
  wire [1:0] filter_0_io_s_axis_tuser_hi = {io_xbar_in_bits_tkeep[14:12] == 3'h4,io_xbar_in_bits_tkeep[10:8] == 3'h4}; // @[BFS.scala 886:106]
  wire  _filter_1_io_s_axis_tkeep_T_3 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[31:0]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_4 = filter_0_m_axis_tkeep[0] & _filter_1_io_s_axis_tkeep_T_3; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_8 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[63:32]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_9 = filter_0_m_axis_tkeep[1] & _filter_1_io_s_axis_tkeep_T_8; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_13 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[95:64]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_14 = filter_0_m_axis_tkeep[2] & _filter_1_io_s_axis_tkeep_T_13; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_18 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[127:96]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_19 = filter_0_m_axis_tkeep[3] & _filter_1_io_s_axis_tkeep_T_18; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_23 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[159:128]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_24 = filter_0_m_axis_tkeep[4] & _filter_1_io_s_axis_tkeep_T_23; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_28 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[191:160]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_29 = filter_0_m_axis_tkeep[5] & _filter_1_io_s_axis_tkeep_T_28; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_33 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[223:192]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_34 = filter_0_m_axis_tkeep[6] & _filter_1_io_s_axis_tkeep_T_33; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_38 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[255:224]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_39 = filter_0_m_axis_tkeep[7] & _filter_1_io_s_axis_tkeep_T_38; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_43 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[287:256]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_44 = filter_0_m_axis_tkeep[8] & _filter_1_io_s_axis_tkeep_T_43; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_48 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[319:288]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_49 = filter_0_m_axis_tkeep[9] & _filter_1_io_s_axis_tkeep_T_48; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_53 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[351:320]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_54 = filter_0_m_axis_tkeep[10] & _filter_1_io_s_axis_tkeep_T_53; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_58 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[383:352]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_59 = filter_0_m_axis_tkeep[11] & _filter_1_io_s_axis_tkeep_T_58; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_63 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[415:384]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_64 = filter_0_m_axis_tkeep[12] & _filter_1_io_s_axis_tkeep_T_63; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_68 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[447:416]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_69 = filter_0_m_axis_tkeep[13] & _filter_1_io_s_axis_tkeep_T_68; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_73 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[479:448]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_74 = filter_0_m_axis_tkeep[14] & _filter_1_io_s_axis_tkeep_T_73; // @[BFS.scala 899:42]
  wire  _filter_1_io_s_axis_tkeep_T_78 = fat_vertex_entry_0_bits[31:0] != filter_0_m_axis_tdata[511:480]; // @[BFS.scala 900:47]
  wire  _filter_1_io_s_axis_tkeep_T_79 = filter_0_m_axis_tkeep[15] & _filter_1_io_s_axis_tkeep_T_78; // @[BFS.scala 899:42]
  wire [7:0] filter_1_io_s_axis_tkeep_lo = {_filter_1_io_s_axis_tkeep_T_39,_filter_1_io_s_axis_tkeep_T_34,
    _filter_1_io_s_axis_tkeep_T_29,_filter_1_io_s_axis_tkeep_T_24,_filter_1_io_s_axis_tkeep_T_19,
    _filter_1_io_s_axis_tkeep_T_14,_filter_1_io_s_axis_tkeep_T_9,_filter_1_io_s_axis_tkeep_T_4}; // @[BFS.scala 902:17]
  wire [15:0] _filter_1_io_s_axis_tkeep_T_80 = {_filter_1_io_s_axis_tkeep_T_79,_filter_1_io_s_axis_tkeep_T_74,
    _filter_1_io_s_axis_tkeep_T_69,_filter_1_io_s_axis_tkeep_T_64,_filter_1_io_s_axis_tkeep_T_59,
    _filter_1_io_s_axis_tkeep_T_54,_filter_1_io_s_axis_tkeep_T_49,_filter_1_io_s_axis_tkeep_T_44,
    filter_1_io_s_axis_tkeep_lo}; // @[BFS.scala 902:17]
  wire  _filter_2_io_s_axis_tkeep_T_3 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[31:0]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_4 = filter_1_m_axis_tkeep[0] & _filter_2_io_s_axis_tkeep_T_3; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_8 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[63:32]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_9 = filter_1_m_axis_tkeep[1] & _filter_2_io_s_axis_tkeep_T_8; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_13 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[95:64]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_14 = filter_1_m_axis_tkeep[2] & _filter_2_io_s_axis_tkeep_T_13; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_18 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[127:96]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_19 = filter_1_m_axis_tkeep[3] & _filter_2_io_s_axis_tkeep_T_18; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_23 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[159:128]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_24 = filter_1_m_axis_tkeep[4] & _filter_2_io_s_axis_tkeep_T_23; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_28 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[191:160]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_29 = filter_1_m_axis_tkeep[5] & _filter_2_io_s_axis_tkeep_T_28; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_33 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[223:192]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_34 = filter_1_m_axis_tkeep[6] & _filter_2_io_s_axis_tkeep_T_33; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_38 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[255:224]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_39 = filter_1_m_axis_tkeep[7] & _filter_2_io_s_axis_tkeep_T_38; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_43 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[287:256]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_44 = filter_1_m_axis_tkeep[8] & _filter_2_io_s_axis_tkeep_T_43; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_48 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[319:288]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_49 = filter_1_m_axis_tkeep[9] & _filter_2_io_s_axis_tkeep_T_48; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_53 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[351:320]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_54 = filter_1_m_axis_tkeep[10] & _filter_2_io_s_axis_tkeep_T_53; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_58 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[383:352]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_59 = filter_1_m_axis_tkeep[11] & _filter_2_io_s_axis_tkeep_T_58; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_63 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[415:384]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_64 = filter_1_m_axis_tkeep[12] & _filter_2_io_s_axis_tkeep_T_63; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_68 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[447:416]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_69 = filter_1_m_axis_tkeep[13] & _filter_2_io_s_axis_tkeep_T_68; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_73 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[479:448]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_74 = filter_1_m_axis_tkeep[14] & _filter_2_io_s_axis_tkeep_T_73; // @[BFS.scala 899:42]
  wire  _filter_2_io_s_axis_tkeep_T_78 = fat_vertex_entry_1_bits[31:0] != filter_1_m_axis_tdata[511:480]; // @[BFS.scala 900:47]
  wire  _filter_2_io_s_axis_tkeep_T_79 = filter_1_m_axis_tkeep[15] & _filter_2_io_s_axis_tkeep_T_78; // @[BFS.scala 899:42]
  wire [7:0] filter_2_io_s_axis_tkeep_lo = {_filter_2_io_s_axis_tkeep_T_39,_filter_2_io_s_axis_tkeep_T_34,
    _filter_2_io_s_axis_tkeep_T_29,_filter_2_io_s_axis_tkeep_T_24,_filter_2_io_s_axis_tkeep_T_19,
    _filter_2_io_s_axis_tkeep_T_14,_filter_2_io_s_axis_tkeep_T_9,_filter_2_io_s_axis_tkeep_T_4}; // @[BFS.scala 902:17]
  wire [15:0] _filter_2_io_s_axis_tkeep_T_80 = {_filter_2_io_s_axis_tkeep_T_79,_filter_2_io_s_axis_tkeep_T_74,
    _filter_2_io_s_axis_tkeep_T_69,_filter_2_io_s_axis_tkeep_T_64,_filter_2_io_s_axis_tkeep_T_59,
    _filter_2_io_s_axis_tkeep_T_54,_filter_2_io_s_axis_tkeep_T_49,_filter_2_io_s_axis_tkeep_T_44,
    filter_2_io_s_axis_tkeep_lo}; // @[BFS.scala 902:17]
  wire  _filter_3_io_s_axis_tkeep_T_3 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[31:0]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_4 = filter_2_m_axis_tkeep[0] & _filter_3_io_s_axis_tkeep_T_3; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_8 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[63:32]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_9 = filter_2_m_axis_tkeep[1] & _filter_3_io_s_axis_tkeep_T_8; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_13 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[95:64]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_14 = filter_2_m_axis_tkeep[2] & _filter_3_io_s_axis_tkeep_T_13; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_18 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[127:96]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_19 = filter_2_m_axis_tkeep[3] & _filter_3_io_s_axis_tkeep_T_18; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_23 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[159:128]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_24 = filter_2_m_axis_tkeep[4] & _filter_3_io_s_axis_tkeep_T_23; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_28 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[191:160]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_29 = filter_2_m_axis_tkeep[5] & _filter_3_io_s_axis_tkeep_T_28; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_33 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[223:192]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_34 = filter_2_m_axis_tkeep[6] & _filter_3_io_s_axis_tkeep_T_33; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_38 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[255:224]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_39 = filter_2_m_axis_tkeep[7] & _filter_3_io_s_axis_tkeep_T_38; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_43 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[287:256]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_44 = filter_2_m_axis_tkeep[8] & _filter_3_io_s_axis_tkeep_T_43; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_48 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[319:288]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_49 = filter_2_m_axis_tkeep[9] & _filter_3_io_s_axis_tkeep_T_48; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_53 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[351:320]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_54 = filter_2_m_axis_tkeep[10] & _filter_3_io_s_axis_tkeep_T_53; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_58 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[383:352]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_59 = filter_2_m_axis_tkeep[11] & _filter_3_io_s_axis_tkeep_T_58; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_63 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[415:384]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_64 = filter_2_m_axis_tkeep[12] & _filter_3_io_s_axis_tkeep_T_63; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_68 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[447:416]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_69 = filter_2_m_axis_tkeep[13] & _filter_3_io_s_axis_tkeep_T_68; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_73 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[479:448]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_74 = filter_2_m_axis_tkeep[14] & _filter_3_io_s_axis_tkeep_T_73; // @[BFS.scala 899:42]
  wire  _filter_3_io_s_axis_tkeep_T_78 = fat_vertex_entry_2_bits[31:0] != filter_2_m_axis_tdata[511:480]; // @[BFS.scala 900:47]
  wire  _filter_3_io_s_axis_tkeep_T_79 = filter_2_m_axis_tkeep[15] & _filter_3_io_s_axis_tkeep_T_78; // @[BFS.scala 899:42]
  wire [7:0] filter_3_io_s_axis_tkeep_lo = {_filter_3_io_s_axis_tkeep_T_39,_filter_3_io_s_axis_tkeep_T_34,
    _filter_3_io_s_axis_tkeep_T_29,_filter_3_io_s_axis_tkeep_T_24,_filter_3_io_s_axis_tkeep_T_19,
    _filter_3_io_s_axis_tkeep_T_14,_filter_3_io_s_axis_tkeep_T_9,_filter_3_io_s_axis_tkeep_T_4}; // @[BFS.scala 902:17]
  wire [15:0] _filter_3_io_s_axis_tkeep_T_80 = {_filter_3_io_s_axis_tkeep_T_79,_filter_3_io_s_axis_tkeep_T_74,
    _filter_3_io_s_axis_tkeep_T_69,_filter_3_io_s_axis_tkeep_T_64,_filter_3_io_s_axis_tkeep_T_59,
    _filter_3_io_s_axis_tkeep_T_54,_filter_3_io_s_axis_tkeep_T_49,_filter_3_io_s_axis_tkeep_T_44,
    filter_3_io_s_axis_tkeep_lo}; // @[BFS.scala 902:17]
  wire  _filter_4_io_s_axis_tkeep_T_3 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[31:0]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_4 = filter_3_m_axis_tkeep[0] & _filter_4_io_s_axis_tkeep_T_3; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_8 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[63:32]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_9 = filter_3_m_axis_tkeep[1] & _filter_4_io_s_axis_tkeep_T_8; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_13 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[95:64]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_14 = filter_3_m_axis_tkeep[2] & _filter_4_io_s_axis_tkeep_T_13; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_18 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[127:96]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_19 = filter_3_m_axis_tkeep[3] & _filter_4_io_s_axis_tkeep_T_18; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_23 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[159:128]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_24 = filter_3_m_axis_tkeep[4] & _filter_4_io_s_axis_tkeep_T_23; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_28 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[191:160]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_29 = filter_3_m_axis_tkeep[5] & _filter_4_io_s_axis_tkeep_T_28; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_33 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[223:192]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_34 = filter_3_m_axis_tkeep[6] & _filter_4_io_s_axis_tkeep_T_33; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_38 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[255:224]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_39 = filter_3_m_axis_tkeep[7] & _filter_4_io_s_axis_tkeep_T_38; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_43 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[287:256]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_44 = filter_3_m_axis_tkeep[8] & _filter_4_io_s_axis_tkeep_T_43; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_48 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[319:288]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_49 = filter_3_m_axis_tkeep[9] & _filter_4_io_s_axis_tkeep_T_48; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_53 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[351:320]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_54 = filter_3_m_axis_tkeep[10] & _filter_4_io_s_axis_tkeep_T_53; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_58 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[383:352]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_59 = filter_3_m_axis_tkeep[11] & _filter_4_io_s_axis_tkeep_T_58; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_63 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[415:384]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_64 = filter_3_m_axis_tkeep[12] & _filter_4_io_s_axis_tkeep_T_63; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_68 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[447:416]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_69 = filter_3_m_axis_tkeep[13] & _filter_4_io_s_axis_tkeep_T_68; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_73 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[479:448]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_74 = filter_3_m_axis_tkeep[14] & _filter_4_io_s_axis_tkeep_T_73; // @[BFS.scala 899:42]
  wire  _filter_4_io_s_axis_tkeep_T_78 = fat_vertex_entry_3_bits[31:0] != filter_3_m_axis_tdata[511:480]; // @[BFS.scala 900:47]
  wire  _filter_4_io_s_axis_tkeep_T_79 = filter_3_m_axis_tkeep[15] & _filter_4_io_s_axis_tkeep_T_78; // @[BFS.scala 899:42]
  wire [7:0] filter_4_io_s_axis_tkeep_lo = {_filter_4_io_s_axis_tkeep_T_39,_filter_4_io_s_axis_tkeep_T_34,
    _filter_4_io_s_axis_tkeep_T_29,_filter_4_io_s_axis_tkeep_T_24,_filter_4_io_s_axis_tkeep_T_19,
    _filter_4_io_s_axis_tkeep_T_14,_filter_4_io_s_axis_tkeep_T_9,_filter_4_io_s_axis_tkeep_T_4}; // @[BFS.scala 902:17]
  wire [15:0] _filter_4_io_s_axis_tkeep_T_80 = {_filter_4_io_s_axis_tkeep_T_79,_filter_4_io_s_axis_tkeep_T_74,
    _filter_4_io_s_axis_tkeep_T_69,_filter_4_io_s_axis_tkeep_T_64,_filter_4_io_s_axis_tkeep_T_59,
    _filter_4_io_s_axis_tkeep_T_54,_filter_4_io_s_axis_tkeep_T_49,_filter_4_io_s_axis_tkeep_T_44,
    filter_4_io_s_axis_tkeep_lo}; // @[BFS.scala 902:17]
  wire [63:0] _io_ddr_out_bits_tkeep_T = filter_4_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  _T_5 = filter_4_m_axis_tvalid & filter_4_m_axis_tready & filter_4_m_axis_tuser[0]; // @[BFS.scala 912:87]
  wire  _T_8 = filter_4_m_axis_tdata[63:32] > fat_vertex_entry_0_bits[63:32]; // @[BFS.scala 914:55]
  wire  _T_9 = _T_5 & _T_8; // @[BFS.scala 913:46]
  wire  _GEN_5 = _T_9 | fat_vertex_entry_0_valid; // @[BFS.scala 914:71 BFS.scala 916:17 BFS.scala 884:46]
  wire  _T_15 = filter_4_m_axis_tvalid & filter_4_m_axis_tready & filter_4_m_axis_tuser[1]; // @[BFS.scala 912:87]
  wire  _T_18 = filter_4_m_axis_tdata[191:160] > fat_vertex_entry_1_bits[63:32]; // @[BFS.scala 914:55]
  wire  _T_19 = _T_15 & _T_18; // @[BFS.scala 913:46]
  wire  _GEN_7 = _T_19 | fat_vertex_entry_1_valid; // @[BFS.scala 914:71 BFS.scala 916:17 BFS.scala 884:46]
  wire  _T_25 = filter_4_m_axis_tvalid & filter_4_m_axis_tready & filter_4_m_axis_tuser[2]; // @[BFS.scala 912:87]
  wire  _T_28 = filter_4_m_axis_tdata[319:288] > fat_vertex_entry_2_bits[63:32]; // @[BFS.scala 914:55]
  wire  _T_29 = _T_25 & _T_28; // @[BFS.scala 913:46]
  wire  _GEN_9 = _T_29 | fat_vertex_entry_2_valid; // @[BFS.scala 914:71 BFS.scala 916:17 BFS.scala 884:46]
  wire  _T_35 = filter_4_m_axis_tvalid & filter_4_m_axis_tready & filter_4_m_axis_tuser[3]; // @[BFS.scala 912:87]
  wire  _T_38 = filter_4_m_axis_tdata[447:416] > fat_vertex_entry_3_bits[63:32]; // @[BFS.scala 914:55]
  wire  _T_39 = _T_35 & _T_38; // @[BFS.scala 913:46]
  wire  _GEN_11 = _T_39 | fat_vertex_entry_3_valid; // @[BFS.scala 914:71 BFS.scala 916:17 BFS.scala 884:46]
  fat_vertex_cache_reg_slice filter_0 ( // @[BFS.scala 882:34]
    .aclk(filter_0_aclk),
    .aresetn(filter_0_aresetn),
    .s_axis_tdata(filter_0_s_axis_tdata),
    .s_axis_tkeep(filter_0_s_axis_tkeep),
    .s_axis_tvalid(filter_0_s_axis_tvalid),
    .s_axis_tready(filter_0_s_axis_tready),
    .s_axis_tlast(filter_0_s_axis_tlast),
    .s_axis_tuser(filter_0_s_axis_tuser),
    .m_axis_tdata(filter_0_m_axis_tdata),
    .m_axis_tkeep(filter_0_m_axis_tkeep),
    .m_axis_tvalid(filter_0_m_axis_tvalid),
    .m_axis_tready(filter_0_m_axis_tready),
    .m_axis_tlast(filter_0_m_axis_tlast),
    .m_axis_tuser(filter_0_m_axis_tuser)
  );
  fat_vertex_cache_reg_slice filter_1 ( // @[BFS.scala 882:34]
    .aclk(filter_1_aclk),
    .aresetn(filter_1_aresetn),
    .s_axis_tdata(filter_1_s_axis_tdata),
    .s_axis_tkeep(filter_1_s_axis_tkeep),
    .s_axis_tvalid(filter_1_s_axis_tvalid),
    .s_axis_tready(filter_1_s_axis_tready),
    .s_axis_tlast(filter_1_s_axis_tlast),
    .s_axis_tuser(filter_1_s_axis_tuser),
    .m_axis_tdata(filter_1_m_axis_tdata),
    .m_axis_tkeep(filter_1_m_axis_tkeep),
    .m_axis_tvalid(filter_1_m_axis_tvalid),
    .m_axis_tready(filter_1_m_axis_tready),
    .m_axis_tlast(filter_1_m_axis_tlast),
    .m_axis_tuser(filter_1_m_axis_tuser)
  );
  fat_vertex_cache_reg_slice filter_2 ( // @[BFS.scala 882:34]
    .aclk(filter_2_aclk),
    .aresetn(filter_2_aresetn),
    .s_axis_tdata(filter_2_s_axis_tdata),
    .s_axis_tkeep(filter_2_s_axis_tkeep),
    .s_axis_tvalid(filter_2_s_axis_tvalid),
    .s_axis_tready(filter_2_s_axis_tready),
    .s_axis_tlast(filter_2_s_axis_tlast),
    .s_axis_tuser(filter_2_s_axis_tuser),
    .m_axis_tdata(filter_2_m_axis_tdata),
    .m_axis_tkeep(filter_2_m_axis_tkeep),
    .m_axis_tvalid(filter_2_m_axis_tvalid),
    .m_axis_tready(filter_2_m_axis_tready),
    .m_axis_tlast(filter_2_m_axis_tlast),
    .m_axis_tuser(filter_2_m_axis_tuser)
  );
  fat_vertex_cache_reg_slice filter_3 ( // @[BFS.scala 882:34]
    .aclk(filter_3_aclk),
    .aresetn(filter_3_aresetn),
    .s_axis_tdata(filter_3_s_axis_tdata),
    .s_axis_tkeep(filter_3_s_axis_tkeep),
    .s_axis_tvalid(filter_3_s_axis_tvalid),
    .s_axis_tready(filter_3_s_axis_tready),
    .s_axis_tlast(filter_3_s_axis_tlast),
    .s_axis_tuser(filter_3_s_axis_tuser),
    .m_axis_tdata(filter_3_m_axis_tdata),
    .m_axis_tkeep(filter_3_m_axis_tkeep),
    .m_axis_tvalid(filter_3_m_axis_tvalid),
    .m_axis_tready(filter_3_m_axis_tready),
    .m_axis_tlast(filter_3_m_axis_tlast),
    .m_axis_tuser(filter_3_m_axis_tuser)
  );
  fat_vertex_cache_reg_slice filter_4 ( // @[BFS.scala 882:34]
    .aclk(filter_4_aclk),
    .aresetn(filter_4_aresetn),
    .s_axis_tdata(filter_4_s_axis_tdata),
    .s_axis_tkeep(filter_4_s_axis_tkeep),
    .s_axis_tvalid(filter_4_s_axis_tvalid),
    .s_axis_tready(filter_4_s_axis_tready),
    .s_axis_tlast(filter_4_s_axis_tlast),
    .s_axis_tuser(filter_4_s_axis_tuser),
    .m_axis_tdata(filter_4_m_axis_tdata),
    .m_axis_tkeep(filter_4_m_axis_tkeep),
    .m_axis_tvalid(filter_4_m_axis_tvalid),
    .m_axis_tready(filter_4_m_axis_tready),
    .m_axis_tlast(filter_4_m_axis_tlast),
    .m_axis_tuser(filter_4_m_axis_tuser)
  );
  assign io_xbar_in_ready = filter_0_s_axis_tready; // @[BFS.scala 887:20]
  assign io_ddr_out_valid = filter_4_m_axis_tvalid; // @[BFS.scala 908:20]
  assign io_ddr_out_bits_tdata = filter_4_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_ddr_out_bits_tkeep = _io_ddr_out_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_ddr_out_bits_tlast = filter_4_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign filter_0_aclk = clock; // @[BFS.scala 889:36]
  assign filter_0_aresetn = ~reset; // @[BFS.scala 890:27]
  assign filter_0_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign filter_0_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign filter_0_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 888:30]
  assign filter_0_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign filter_0_s_axis_tuser = {filter_0_io_s_axis_tuser_hi,filter_0_io_s_axis_tuser_lo}; // @[BFS.scala 886:106]
  assign filter_0_m_axis_tready = filter_1_s_axis_tready; // @[BFS.scala 895:19]
  assign filter_1_aclk = clock; // @[BFS.scala 893:32]
  assign filter_1_aresetn = ~reset; // @[BFS.scala 894:23]
  assign filter_1_s_axis_tdata = filter_0_m_axis_tdata; // @[BFS.scala 895:19]
  assign filter_1_s_axis_tkeep = fat_vertex_entry_0_valid ? {{48'd0}, _filter_1_io_s_axis_tkeep_T_80} :
    filter_0_m_axis_tkeep; // @[BFS.scala 896:38 BFS.scala 897:27 BFS.scala 895:19]
  assign filter_1_s_axis_tvalid = filter_0_m_axis_tvalid; // @[BFS.scala 895:19]
  assign filter_1_s_axis_tlast = filter_0_m_axis_tlast; // @[BFS.scala 895:19]
  assign filter_1_s_axis_tuser = filter_0_m_axis_tuser; // @[BFS.scala 895:19]
  assign filter_1_m_axis_tready = filter_2_s_axis_tready; // @[BFS.scala 895:19]
  assign filter_2_aclk = clock; // @[BFS.scala 893:32]
  assign filter_2_aresetn = ~reset; // @[BFS.scala 894:23]
  assign filter_2_s_axis_tdata = filter_1_m_axis_tdata; // @[BFS.scala 895:19]
  assign filter_2_s_axis_tkeep = fat_vertex_entry_1_valid ? {{48'd0}, _filter_2_io_s_axis_tkeep_T_80} :
    filter_1_m_axis_tkeep; // @[BFS.scala 896:38 BFS.scala 897:27 BFS.scala 895:19]
  assign filter_2_s_axis_tvalid = filter_1_m_axis_tvalid; // @[BFS.scala 895:19]
  assign filter_2_s_axis_tlast = filter_1_m_axis_tlast; // @[BFS.scala 895:19]
  assign filter_2_s_axis_tuser = filter_1_m_axis_tuser; // @[BFS.scala 895:19]
  assign filter_2_m_axis_tready = filter_3_s_axis_tready; // @[BFS.scala 895:19]
  assign filter_3_aclk = clock; // @[BFS.scala 893:32]
  assign filter_3_aresetn = ~reset; // @[BFS.scala 894:23]
  assign filter_3_s_axis_tdata = filter_2_m_axis_tdata; // @[BFS.scala 895:19]
  assign filter_3_s_axis_tkeep = fat_vertex_entry_2_valid ? {{48'd0}, _filter_3_io_s_axis_tkeep_T_80} :
    filter_2_m_axis_tkeep; // @[BFS.scala 896:38 BFS.scala 897:27 BFS.scala 895:19]
  assign filter_3_s_axis_tvalid = filter_2_m_axis_tvalid; // @[BFS.scala 895:19]
  assign filter_3_s_axis_tlast = filter_2_m_axis_tlast; // @[BFS.scala 895:19]
  assign filter_3_s_axis_tuser = filter_2_m_axis_tuser; // @[BFS.scala 895:19]
  assign filter_3_m_axis_tready = filter_4_s_axis_tready; // @[BFS.scala 895:19]
  assign filter_4_aclk = clock; // @[BFS.scala 893:32]
  assign filter_4_aresetn = ~reset; // @[BFS.scala 894:23]
  assign filter_4_s_axis_tdata = filter_3_m_axis_tdata; // @[BFS.scala 895:19]
  assign filter_4_s_axis_tkeep = fat_vertex_entry_3_valid ? {{48'd0}, _filter_4_io_s_axis_tkeep_T_80} :
    filter_3_m_axis_tkeep; // @[BFS.scala 896:38 BFS.scala 897:27 BFS.scala 895:19]
  assign filter_4_s_axis_tvalid = filter_3_m_axis_tvalid; // @[BFS.scala 895:19]
  assign filter_4_s_axis_tlast = filter_3_m_axis_tlast; // @[BFS.scala 895:19]
  assign filter_4_s_axis_tuser = filter_3_m_axis_tuser; // @[BFS.scala 895:19]
  assign filter_4_m_axis_tready = io_ddr_out_ready; // @[BFS.scala 907:30]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 884:46]
      fat_vertex_entry_0_valid <= 1'h0; // @[BFS.scala 884:46]
    end else begin
      fat_vertex_entry_0_valid <= _GEN_5;
    end
    if (reset) begin // @[BFS.scala 884:46]
      fat_vertex_entry_0_bits <= 64'h0; // @[BFS.scala 884:46]
    end else if (_T_9) begin // @[BFS.scala 914:71]
      fat_vertex_entry_0_bits <= filter_4_m_axis_tdata[63:0]; // @[BFS.scala 915:16]
    end
    if (reset) begin // @[BFS.scala 884:46]
      fat_vertex_entry_1_valid <= 1'h0; // @[BFS.scala 884:46]
    end else begin
      fat_vertex_entry_1_valid <= _GEN_7;
    end
    if (reset) begin // @[BFS.scala 884:46]
      fat_vertex_entry_1_bits <= 64'h0; // @[BFS.scala 884:46]
    end else if (_T_19) begin // @[BFS.scala 914:71]
      fat_vertex_entry_1_bits <= filter_4_m_axis_tdata[191:128]; // @[BFS.scala 915:16]
    end
    if (reset) begin // @[BFS.scala 884:46]
      fat_vertex_entry_2_valid <= 1'h0; // @[BFS.scala 884:46]
    end else begin
      fat_vertex_entry_2_valid <= _GEN_9;
    end
    if (reset) begin // @[BFS.scala 884:46]
      fat_vertex_entry_2_bits <= 64'h0; // @[BFS.scala 884:46]
    end else if (_T_29) begin // @[BFS.scala 914:71]
      fat_vertex_entry_2_bits <= filter_4_m_axis_tdata[319:256]; // @[BFS.scala 915:16]
    end
    if (reset) begin // @[BFS.scala 884:46]
      fat_vertex_entry_3_valid <= 1'h0; // @[BFS.scala 884:46]
    end else begin
      fat_vertex_entry_3_valid <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 884:46]
      fat_vertex_entry_3_bits <= 64'h0; // @[BFS.scala 884:46]
    end else if (_T_39) begin // @[BFS.scala 914:71]
      fat_vertex_entry_3_bits <= filter_4_m_axis_tdata[447:384]; // @[BFS.scala 915:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fat_vertex_entry_0_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  fat_vertex_entry_0_bits = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  fat_vertex_entry_1_valid = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  fat_vertex_entry_1_bits = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  fat_vertex_entry_2_valid = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  fat_vertex_entry_2_bits = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  fat_vertex_entry_3_valid = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  fat_vertex_entry_3_bits = _RAND_7[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module broadcast_xbar(
  input          clock,
  input          reset,
  output         io_ddr_in_0_ready,
  input          io_ddr_in_0_valid,
  input  [127:0] io_ddr_in_0_bits_tdata,
  input  [3:0]   io_ddr_in_0_bits_tkeep,
  input          io_ddr_in_0_bits_tlast,
  output         io_ddr_in_1_ready,
  input          io_ddr_in_1_valid,
  input  [127:0] io_ddr_in_1_bits_tdata,
  input  [3:0]   io_ddr_in_1_bits_tkeep,
  input          io_ddr_in_1_bits_tlast,
  output         io_ddr_in_2_ready,
  input          io_ddr_in_2_valid,
  input  [127:0] io_ddr_in_2_bits_tdata,
  input  [3:0]   io_ddr_in_2_bits_tkeep,
  input          io_ddr_in_2_bits_tlast,
  output         io_ddr_in_3_ready,
  input          io_ddr_in_3_valid,
  input  [127:0] io_ddr_in_3_bits_tdata,
  input  [3:0]   io_ddr_in_3_bits_tkeep,
  input          io_ddr_in_3_bits_tlast,
  input          io_pe_out_0_ready,
  output         io_pe_out_0_valid,
  output [511:0] io_pe_out_0_bits_tdata,
  output [15:0]  io_pe_out_0_bits_tkeep,
  output         io_pe_out_0_bits_tlast,
  input          io_pe_out_1_ready,
  output         io_pe_out_1_valid,
  output [511:0] io_pe_out_1_bits_tdata,
  output [15:0]  io_pe_out_1_bits_tkeep,
  output         io_pe_out_1_bits_tlast,
  input          io_pe_out_2_ready,
  output         io_pe_out_2_valid,
  output [511:0] io_pe_out_2_bits_tdata,
  output [15:0]  io_pe_out_2_bits_tkeep,
  output         io_pe_out_2_bits_tlast,
  input          io_pe_out_3_ready,
  output         io_pe_out_3_valid,
  output [511:0] io_pe_out_3_bits_tdata,
  output [15:0]  io_pe_out_3_bits_tkeep,
  output         io_pe_out_3_bits_tlast,
  input          io_pe_out_4_ready,
  output         io_pe_out_4_valid,
  output [511:0] io_pe_out_4_bits_tdata,
  output [15:0]  io_pe_out_4_bits_tkeep,
  output         io_pe_out_4_bits_tlast,
  input          io_pe_out_5_ready,
  output         io_pe_out_5_valid,
  output [511:0] io_pe_out_5_bits_tdata,
  output [15:0]  io_pe_out_5_bits_tkeep,
  output         io_pe_out_5_bits_tlast,
  input          io_pe_out_6_ready,
  output         io_pe_out_6_valid,
  output [511:0] io_pe_out_6_bits_tdata,
  output [15:0]  io_pe_out_6_bits_tkeep,
  output         io_pe_out_6_bits_tlast,
  input          io_pe_out_7_ready,
  output         io_pe_out_7_valid,
  output [511:0] io_pe_out_7_bits_tdata,
  output [15:0]  io_pe_out_7_bits_tkeep,
  output         io_pe_out_7_bits_tlast,
  input          io_pe_out_8_ready,
  output         io_pe_out_8_valid,
  output [511:0] io_pe_out_8_bits_tdata,
  output [15:0]  io_pe_out_8_bits_tkeep,
  output         io_pe_out_8_bits_tlast,
  input          io_pe_out_9_ready,
  output         io_pe_out_9_valid,
  output [511:0] io_pe_out_9_bits_tdata,
  output [15:0]  io_pe_out_9_bits_tkeep,
  output         io_pe_out_9_bits_tlast,
  input          io_pe_out_10_ready,
  output         io_pe_out_10_valid,
  output [511:0] io_pe_out_10_bits_tdata,
  output [15:0]  io_pe_out_10_bits_tkeep,
  output         io_pe_out_10_bits_tlast,
  input          io_pe_out_11_ready,
  output         io_pe_out_11_valid,
  output [511:0] io_pe_out_11_bits_tdata,
  output [15:0]  io_pe_out_11_bits_tkeep,
  output         io_pe_out_11_bits_tlast,
  input          io_pe_out_12_ready,
  output         io_pe_out_12_valid,
  output [511:0] io_pe_out_12_bits_tdata,
  output [15:0]  io_pe_out_12_bits_tkeep,
  output         io_pe_out_12_bits_tlast,
  input          io_pe_out_13_ready,
  output         io_pe_out_13_valid,
  output [511:0] io_pe_out_13_bits_tdata,
  output [15:0]  io_pe_out_13_bits_tkeep,
  output         io_pe_out_13_bits_tlast,
  input          io_pe_out_14_ready,
  output         io_pe_out_14_valid,
  output [511:0] io_pe_out_14_bits_tdata,
  output [15:0]  io_pe_out_14_bits_tkeep,
  output         io_pe_out_14_bits_tlast,
  input          io_pe_out_15_ready,
  output         io_pe_out_15_valid,
  output [511:0] io_pe_out_15_bits_tdata,
  output [15:0]  io_pe_out_15_bits_tkeep,
  output         io_pe_out_15_bits_tlast
);
  wire  xbar_aclk; // @[BFS.scala 931:20]
  wire  xbar_aresetn; // @[BFS.scala 931:20]
  wire [511:0] xbar_s_axis_tdata; // @[BFS.scala 931:20]
  wire [63:0] xbar_s_axis_tkeep; // @[BFS.scala 931:20]
  wire  xbar_s_axis_tvalid; // @[BFS.scala 931:20]
  wire  xbar_s_axis_tready; // @[BFS.scala 931:20]
  wire  xbar_s_axis_tlast; // @[BFS.scala 931:20]
  wire  xbar_s_axis_tid; // @[BFS.scala 931:20]
  wire [8191:0] xbar_m_axis_tdata; // @[BFS.scala 931:20]
  wire [1023:0] xbar_m_axis_tkeep; // @[BFS.scala 931:20]
  wire [15:0] xbar_m_axis_tvalid; // @[BFS.scala 931:20]
  wire [15:0] xbar_m_axis_tready; // @[BFS.scala 931:20]
  wire [15:0] xbar_m_axis_tlast; // @[BFS.scala 931:20]
  wire [15:0] xbar_m_axis_tid; // @[BFS.scala 931:20]
  wire  combiner_aclk; // @[BFS.scala 938:26]
  wire  combiner_aresetn; // @[BFS.scala 938:26]
  wire [511:0] combiner_s_axis_tdata; // @[BFS.scala 938:26]
  wire [63:0] combiner_s_axis_tkeep; // @[BFS.scala 938:26]
  wire [3:0] combiner_s_axis_tvalid; // @[BFS.scala 938:26]
  wire [3:0] combiner_s_axis_tready; // @[BFS.scala 938:26]
  wire [3:0] combiner_s_axis_tlast; // @[BFS.scala 938:26]
  wire [3:0] combiner_s_axis_tid; // @[BFS.scala 938:26]
  wire [511:0] combiner_m_axis_tdata; // @[BFS.scala 938:26]
  wire [63:0] combiner_m_axis_tkeep; // @[BFS.scala 938:26]
  wire  combiner_m_axis_tvalid; // @[BFS.scala 938:26]
  wire  combiner_m_axis_tready; // @[BFS.scala 938:26]
  wire  combiner_m_axis_tlast; // @[BFS.scala 938:26]
  wire  combiner_m_axis_tid; // @[BFS.scala 938:26]
  wire  buffer0_s_axis_aclk; // @[BFS.scala 950:25]
  wire  buffer0_s_axis_aresetn; // @[BFS.scala 950:25]
  wire [511:0] buffer0_s_axis_tdata; // @[BFS.scala 950:25]
  wire [63:0] buffer0_s_axis_tkeep; // @[BFS.scala 950:25]
  wire  buffer0_s_axis_tvalid; // @[BFS.scala 950:25]
  wire  buffer0_s_axis_tready; // @[BFS.scala 950:25]
  wire  buffer0_s_axis_tlast; // @[BFS.scala 950:25]
  wire  buffer0_s_axis_tid; // @[BFS.scala 950:25]
  wire [511:0] buffer0_m_axis_tdata; // @[BFS.scala 950:25]
  wire [63:0] buffer0_m_axis_tkeep; // @[BFS.scala 950:25]
  wire  buffer0_m_axis_tvalid; // @[BFS.scala 950:25]
  wire  buffer0_m_axis_tready; // @[BFS.scala 950:25]
  wire  buffer0_m_axis_tlast; // @[BFS.scala 950:25]
  wire  buffer0_m_axis_tid; // @[BFS.scala 950:25]
  wire  fat_vertex_filter_clock; // @[BFS.scala 955:35]
  wire  fat_vertex_filter_reset; // @[BFS.scala 955:35]
  wire  fat_vertex_filter_io_xbar_in_ready; // @[BFS.scala 955:35]
  wire  fat_vertex_filter_io_xbar_in_valid; // @[BFS.scala 955:35]
  wire [511:0] fat_vertex_filter_io_xbar_in_bits_tdata; // @[BFS.scala 955:35]
  wire [15:0] fat_vertex_filter_io_xbar_in_bits_tkeep; // @[BFS.scala 955:35]
  wire  fat_vertex_filter_io_xbar_in_bits_tlast; // @[BFS.scala 955:35]
  wire  fat_vertex_filter_io_ddr_out_ready; // @[BFS.scala 955:35]
  wire  fat_vertex_filter_io_ddr_out_valid; // @[BFS.scala 955:35]
  wire [511:0] fat_vertex_filter_io_ddr_out_bits_tdata; // @[BFS.scala 955:35]
  wire [15:0] fat_vertex_filter_io_ddr_out_bits_tkeep; // @[BFS.scala 955:35]
  wire  fat_vertex_filter_io_ddr_out_bits_tlast; // @[BFS.scala 955:35]
  wire [255:0] combiner_io_s_axis_tdata_lo = {io_ddr_in_1_bits_tdata,io_ddr_in_0_bits_tdata}; // @[BFS.scala 941:98]
  wire [255:0] combiner_io_s_axis_tdata_hi = {io_ddr_in_3_bits_tdata,io_ddr_in_2_bits_tdata}; // @[BFS.scala 941:98]
  wire  _combiner_io_s_axis_tkeep_T_4 = io_ddr_in_0_bits_tkeep[0] & io_ddr_in_0_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_5 = io_ddr_in_0_bits_tkeep[1] & io_ddr_in_0_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_6 = io_ddr_in_0_bits_tkeep[2] & io_ddr_in_0_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_7 = io_ddr_in_0_bits_tkeep[3] & io_ddr_in_0_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_12 = io_ddr_in_1_bits_tkeep[0] & io_ddr_in_1_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_13 = io_ddr_in_1_bits_tkeep[1] & io_ddr_in_1_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_14 = io_ddr_in_1_bits_tkeep[2] & io_ddr_in_1_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_15 = io_ddr_in_1_bits_tkeep[3] & io_ddr_in_1_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_20 = io_ddr_in_2_bits_tkeep[0] & io_ddr_in_2_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_21 = io_ddr_in_2_bits_tkeep[1] & io_ddr_in_2_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_22 = io_ddr_in_2_bits_tkeep[2] & io_ddr_in_2_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_23 = io_ddr_in_2_bits_tkeep[3] & io_ddr_in_2_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_28 = io_ddr_in_3_bits_tkeep[0] & io_ddr_in_3_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_29 = io_ddr_in_3_bits_tkeep[1] & io_ddr_in_3_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_30 = io_ddr_in_3_bits_tkeep[2] & io_ddr_in_3_valid; // @[BFS.scala 942:120]
  wire  _combiner_io_s_axis_tkeep_T_31 = io_ddr_in_3_bits_tkeep[3] & io_ddr_in_3_valid; // @[BFS.scala 942:120]
  wire [7:0] combiner_io_s_axis_tkeep_lo = {_combiner_io_s_axis_tkeep_T_15,_combiner_io_s_axis_tkeep_T_14,
    _combiner_io_s_axis_tkeep_T_13,_combiner_io_s_axis_tkeep_T_12,_combiner_io_s_axis_tkeep_T_7,
    _combiner_io_s_axis_tkeep_T_6,_combiner_io_s_axis_tkeep_T_5,_combiner_io_s_axis_tkeep_T_4}; // @[BFS.scala 943:35]
  wire [15:0] _combiner_io_s_axis_tkeep_T_32 = {_combiner_io_s_axis_tkeep_T_31,_combiner_io_s_axis_tkeep_T_30,
    _combiner_io_s_axis_tkeep_T_29,_combiner_io_s_axis_tkeep_T_28,_combiner_io_s_axis_tkeep_T_23,
    _combiner_io_s_axis_tkeep_T_22,_combiner_io_s_axis_tkeep_T_21,_combiner_io_s_axis_tkeep_T_20,
    combiner_io_s_axis_tkeep_lo}; // @[BFS.scala 943:35]
  wire [1:0] combiner_io_s_axis_tlast_lo = {io_ddr_in_1_bits_tlast,io_ddr_in_0_bits_tlast}; // @[BFS.scala 944:98]
  wire [1:0] combiner_io_s_axis_tlast_hi = {io_ddr_in_3_bits_tlast,io_ddr_in_2_bits_tlast}; // @[BFS.scala 944:98]
  wire  _combiner_io_s_axis_tvalid_T_2 = io_ddr_in_0_valid | io_ddr_in_1_valid | io_ddr_in_2_valid | io_ddr_in_3_valid; // @[BFS.scala 945:99]
  wire [1:0] combiner_io_s_axis_tvalid_lo = {_combiner_io_s_axis_tvalid_T_2,_combiner_io_s_axis_tvalid_T_2}; // @[BFS.scala 945:111]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_64 = buffer0_m_axis_tkeep[0] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_65 = buffer0_m_axis_tkeep[1] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_66 = buffer0_m_axis_tkeep[2] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_67 = buffer0_m_axis_tkeep[3] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_68 = buffer0_m_axis_tkeep[4] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_69 = buffer0_m_axis_tkeep[5] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_70 = buffer0_m_axis_tkeep[6] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_71 = buffer0_m_axis_tkeep[7] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_72 = buffer0_m_axis_tkeep[8] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_73 = buffer0_m_axis_tkeep[9] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_74 = buffer0_m_axis_tkeep[10] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_75 = buffer0_m_axis_tkeep[11] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_76 = buffer0_m_axis_tkeep[12] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_77 = buffer0_m_axis_tkeep[13] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_78 = buffer0_m_axis_tkeep[14] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_79 = buffer0_m_axis_tkeep[15] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_80 = buffer0_m_axis_tkeep[16] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_81 = buffer0_m_axis_tkeep[17] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_82 = buffer0_m_axis_tkeep[18] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_83 = buffer0_m_axis_tkeep[19] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_84 = buffer0_m_axis_tkeep[20] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_85 = buffer0_m_axis_tkeep[21] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_86 = buffer0_m_axis_tkeep[22] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_87 = buffer0_m_axis_tkeep[23] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_88 = buffer0_m_axis_tkeep[24] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_89 = buffer0_m_axis_tkeep[25] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_90 = buffer0_m_axis_tkeep[26] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_91 = buffer0_m_axis_tkeep[27] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_92 = buffer0_m_axis_tkeep[28] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_93 = buffer0_m_axis_tkeep[29] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_94 = buffer0_m_axis_tkeep[30] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_95 = buffer0_m_axis_tkeep[31] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_96 = buffer0_m_axis_tkeep[32] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_97 = buffer0_m_axis_tkeep[33] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_98 = buffer0_m_axis_tkeep[34] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_99 = buffer0_m_axis_tkeep[35] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_100 = buffer0_m_axis_tkeep[36] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_101 = buffer0_m_axis_tkeep[37] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_102 = buffer0_m_axis_tkeep[38] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_103 = buffer0_m_axis_tkeep[39] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_104 = buffer0_m_axis_tkeep[40] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_105 = buffer0_m_axis_tkeep[41] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_106 = buffer0_m_axis_tkeep[42] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_107 = buffer0_m_axis_tkeep[43] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_108 = buffer0_m_axis_tkeep[44] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_109 = buffer0_m_axis_tkeep[45] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_110 = buffer0_m_axis_tkeep[46] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_111 = buffer0_m_axis_tkeep[47] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_112 = buffer0_m_axis_tkeep[48] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_113 = buffer0_m_axis_tkeep[49] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_114 = buffer0_m_axis_tkeep[50] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_115 = buffer0_m_axis_tkeep[51] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_116 = buffer0_m_axis_tkeep[52] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_117 = buffer0_m_axis_tkeep[53] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_118 = buffer0_m_axis_tkeep[54] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_119 = buffer0_m_axis_tkeep[55] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_120 = buffer0_m_axis_tkeep[56] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_121 = buffer0_m_axis_tkeep[57] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_122 = buffer0_m_axis_tkeep[58] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_123 = buffer0_m_axis_tkeep[59] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_124 = buffer0_m_axis_tkeep[60] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_125 = buffer0_m_axis_tkeep[61] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_126 = buffer0_m_axis_tkeep[62] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire  _fat_vertex_filter_io_xbar_in_bits_tkeep_T_127 = buffer0_m_axis_tkeep[63] & buffer0_m_axis_tvalid; // @[BFS.scala 958:60]
  wire [7:0] fat_vertex_filter_io_xbar_in_bits_tkeep_lo_lo_lo = {_fat_vertex_filter_io_xbar_in_bits_tkeep_T_71,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_70,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_69,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_68,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_67,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_66,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_65,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_64}; // @[BFS.scala 958:95]
  wire [15:0] fat_vertex_filter_io_xbar_in_bits_tkeep_lo_lo = {_fat_vertex_filter_io_xbar_in_bits_tkeep_T_79,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_78,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_77,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_76,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_75,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_74,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_73,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_72,fat_vertex_filter_io_xbar_in_bits_tkeep_lo_lo_lo}; // @[BFS.scala 958:95]
  wire [7:0] fat_vertex_filter_io_xbar_in_bits_tkeep_lo_hi_lo = {_fat_vertex_filter_io_xbar_in_bits_tkeep_T_87,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_86,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_85,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_84,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_83,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_82,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_81,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_80}; // @[BFS.scala 958:95]
  wire [31:0] fat_vertex_filter_io_xbar_in_bits_tkeep_lo = {_fat_vertex_filter_io_xbar_in_bits_tkeep_T_95,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_94,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_93,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_92,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_91,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_90,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_89,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_88,fat_vertex_filter_io_xbar_in_bits_tkeep_lo_hi_lo,
    fat_vertex_filter_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 958:95]
  wire [7:0] fat_vertex_filter_io_xbar_in_bits_tkeep_hi_lo_lo = {_fat_vertex_filter_io_xbar_in_bits_tkeep_T_103,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_102,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_101,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_100,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_99,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_98,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_97,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_96}; // @[BFS.scala 958:95]
  wire [15:0] fat_vertex_filter_io_xbar_in_bits_tkeep_hi_lo = {_fat_vertex_filter_io_xbar_in_bits_tkeep_T_111,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_110,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_109,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_108,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_107,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_106,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_105,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_104,fat_vertex_filter_io_xbar_in_bits_tkeep_hi_lo_lo}; // @[BFS.scala 958:95]
  wire [7:0] fat_vertex_filter_io_xbar_in_bits_tkeep_hi_hi_lo = {_fat_vertex_filter_io_xbar_in_bits_tkeep_T_119,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_118,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_117,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_116,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_115,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_114,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_113,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_112}; // @[BFS.scala 958:95]
  wire [31:0] fat_vertex_filter_io_xbar_in_bits_tkeep_hi = {_fat_vertex_filter_io_xbar_in_bits_tkeep_T_127,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_126,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_125,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_124,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_123,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_122,_fat_vertex_filter_io_xbar_in_bits_tkeep_T_121,
    _fat_vertex_filter_io_xbar_in_bits_tkeep_T_120,fat_vertex_filter_io_xbar_in_bits_tkeep_hi_hi_lo,
    fat_vertex_filter_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 958:95]
  wire [63:0] _fat_vertex_filter_io_xbar_in_bits_tkeep_T_128 = {fat_vertex_filter_io_xbar_in_bits_tkeep_hi,
    fat_vertex_filter_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 958:95]
  wire [7:0] xbar_io_m_axis_tready_lo = {io_pe_out_7_ready,io_pe_out_6_ready,io_pe_out_5_ready,io_pe_out_4_ready,
    io_pe_out_3_ready,io_pe_out_2_ready,io_pe_out_1_ready,io_pe_out_0_ready}; // @[BFS.scala 978:12]
  wire [7:0] xbar_io_m_axis_tready_hi = {io_pe_out_15_ready,io_pe_out_14_ready,io_pe_out_13_ready,io_pe_out_12_ready,
    io_pe_out_11_ready,io_pe_out_10_ready,io_pe_out_9_ready,io_pe_out_8_ready}; // @[BFS.scala 978:12]
  axis_broadcaster_64 xbar ( // @[BFS.scala 931:20]
    .aclk(xbar_aclk),
    .aresetn(xbar_aresetn),
    .s_axis_tdata(xbar_s_axis_tdata),
    .s_axis_tkeep(xbar_s_axis_tkeep),
    .s_axis_tvalid(xbar_s_axis_tvalid),
    .s_axis_tready(xbar_s_axis_tready),
    .s_axis_tlast(xbar_s_axis_tlast),
    .s_axis_tid(xbar_s_axis_tid),
    .m_axis_tdata(xbar_m_axis_tdata),
    .m_axis_tkeep(xbar_m_axis_tkeep),
    .m_axis_tvalid(xbar_m_axis_tvalid),
    .m_axis_tready(xbar_m_axis_tready),
    .m_axis_tlast(xbar_m_axis_tlast),
    .m_axis_tid(xbar_m_axis_tid)
  );
  axis_combiner_level0 combiner ( // @[BFS.scala 938:26]
    .aclk(combiner_aclk),
    .aresetn(combiner_aresetn),
    .s_axis_tdata(combiner_s_axis_tdata),
    .s_axis_tkeep(combiner_s_axis_tkeep),
    .s_axis_tvalid(combiner_s_axis_tvalid),
    .s_axis_tready(combiner_s_axis_tready),
    .s_axis_tlast(combiner_s_axis_tlast),
    .s_axis_tid(combiner_s_axis_tid),
    .m_axis_tdata(combiner_m_axis_tdata),
    .m_axis_tkeep(combiner_m_axis_tkeep),
    .m_axis_tvalid(combiner_m_axis_tvalid),
    .m_axis_tready(combiner_m_axis_tready),
    .m_axis_tlast(combiner_m_axis_tlast),
    .m_axis_tid(combiner_m_axis_tid)
  );
  Remote_xbar_buffer0 buffer0 ( // @[BFS.scala 950:25]
    .s_axis_aclk(buffer0_s_axis_aclk),
    .s_axis_aresetn(buffer0_s_axis_aresetn),
    .s_axis_tdata(buffer0_s_axis_tdata),
    .s_axis_tkeep(buffer0_s_axis_tkeep),
    .s_axis_tvalid(buffer0_s_axis_tvalid),
    .s_axis_tready(buffer0_s_axis_tready),
    .s_axis_tlast(buffer0_s_axis_tlast),
    .s_axis_tid(buffer0_s_axis_tid),
    .m_axis_tdata(buffer0_m_axis_tdata),
    .m_axis_tkeep(buffer0_m_axis_tkeep),
    .m_axis_tvalid(buffer0_m_axis_tvalid),
    .m_axis_tready(buffer0_m_axis_tready),
    .m_axis_tlast(buffer0_m_axis_tlast),
    .m_axis_tid(buffer0_m_axis_tid)
  );
  fat_vertex_cache fat_vertex_filter ( // @[BFS.scala 955:35]
    .clock(fat_vertex_filter_clock),
    .reset(fat_vertex_filter_reset),
    .io_xbar_in_ready(fat_vertex_filter_io_xbar_in_ready),
    .io_xbar_in_valid(fat_vertex_filter_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(fat_vertex_filter_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(fat_vertex_filter_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(fat_vertex_filter_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(fat_vertex_filter_io_ddr_out_ready),
    .io_ddr_out_valid(fat_vertex_filter_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(fat_vertex_filter_io_ddr_out_bits_tdata),
    .io_ddr_out_bits_tkeep(fat_vertex_filter_io_ddr_out_bits_tkeep),
    .io_ddr_out_bits_tlast(fat_vertex_filter_io_ddr_out_bits_tlast)
  );
  assign io_ddr_in_0_ready = combiner_s_axis_tready[0]; // @[BFS.scala 947:60]
  assign io_ddr_in_1_ready = combiner_s_axis_tready[1]; // @[BFS.scala 947:60]
  assign io_ddr_in_2_ready = combiner_s_axis_tready[2]; // @[BFS.scala 947:60]
  assign io_ddr_in_3_ready = combiner_s_axis_tready[3]; // @[BFS.scala 947:60]
  assign io_pe_out_0_valid = xbar_m_axis_tvalid[0]; // @[BFS.scala 973:40]
  assign io_pe_out_0_bits_tdata = xbar_m_axis_tdata[511:0]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_0_bits_tkeep = xbar_m_axis_tkeep[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_0_bits_tlast = xbar_m_axis_tlast[0]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_1_valid = xbar_m_axis_tvalid[1]; // @[BFS.scala 973:40]
  assign io_pe_out_1_bits_tdata = xbar_m_axis_tdata[1023:512]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_1_bits_tkeep = xbar_m_axis_tkeep[79:64]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_1_bits_tlast = xbar_m_axis_tlast[1]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_2_valid = xbar_m_axis_tvalid[2]; // @[BFS.scala 973:40]
  assign io_pe_out_2_bits_tdata = xbar_m_axis_tdata[1535:1024]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_2_bits_tkeep = xbar_m_axis_tkeep[143:128]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_2_bits_tlast = xbar_m_axis_tlast[2]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_3_valid = xbar_m_axis_tvalid[3]; // @[BFS.scala 973:40]
  assign io_pe_out_3_bits_tdata = xbar_m_axis_tdata[2047:1536]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_3_bits_tkeep = xbar_m_axis_tkeep[207:192]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_3_bits_tlast = xbar_m_axis_tlast[3]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_4_valid = xbar_m_axis_tvalid[4]; // @[BFS.scala 973:40]
  assign io_pe_out_4_bits_tdata = xbar_m_axis_tdata[2559:2048]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_4_bits_tkeep = xbar_m_axis_tkeep[271:256]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_4_bits_tlast = xbar_m_axis_tlast[4]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_5_valid = xbar_m_axis_tvalid[5]; // @[BFS.scala 973:40]
  assign io_pe_out_5_bits_tdata = xbar_m_axis_tdata[3071:2560]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_5_bits_tkeep = xbar_m_axis_tkeep[335:320]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_5_bits_tlast = xbar_m_axis_tlast[5]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_6_valid = xbar_m_axis_tvalid[6]; // @[BFS.scala 973:40]
  assign io_pe_out_6_bits_tdata = xbar_m_axis_tdata[3583:3072]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_6_bits_tkeep = xbar_m_axis_tkeep[399:384]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_6_bits_tlast = xbar_m_axis_tlast[6]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_7_valid = xbar_m_axis_tvalid[7]; // @[BFS.scala 973:40]
  assign io_pe_out_7_bits_tdata = xbar_m_axis_tdata[4095:3584]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_7_bits_tkeep = xbar_m_axis_tkeep[463:448]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_7_bits_tlast = xbar_m_axis_tlast[7]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_8_valid = xbar_m_axis_tvalid[8]; // @[BFS.scala 973:40]
  assign io_pe_out_8_bits_tdata = xbar_m_axis_tdata[4607:4096]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_8_bits_tkeep = xbar_m_axis_tkeep[527:512]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_8_bits_tlast = xbar_m_axis_tlast[8]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_9_valid = xbar_m_axis_tvalid[9]; // @[BFS.scala 973:40]
  assign io_pe_out_9_bits_tdata = xbar_m_axis_tdata[5119:4608]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_9_bits_tkeep = xbar_m_axis_tkeep[591:576]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_9_bits_tlast = xbar_m_axis_tlast[9]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_10_valid = xbar_m_axis_tvalid[10]; // @[BFS.scala 973:40]
  assign io_pe_out_10_bits_tdata = xbar_m_axis_tdata[5631:5120]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_10_bits_tkeep = xbar_m_axis_tkeep[655:640]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_10_bits_tlast = xbar_m_axis_tlast[10]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_11_valid = xbar_m_axis_tvalid[11]; // @[BFS.scala 973:40]
  assign io_pe_out_11_bits_tdata = xbar_m_axis_tdata[6143:5632]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_11_bits_tkeep = xbar_m_axis_tkeep[719:704]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_11_bits_tlast = xbar_m_axis_tlast[11]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_12_valid = xbar_m_axis_tvalid[12]; // @[BFS.scala 973:40]
  assign io_pe_out_12_bits_tdata = xbar_m_axis_tdata[6655:6144]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_12_bits_tkeep = xbar_m_axis_tkeep[783:768]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_12_bits_tlast = xbar_m_axis_tlast[12]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_13_valid = xbar_m_axis_tvalid[13]; // @[BFS.scala 973:40]
  assign io_pe_out_13_bits_tdata = xbar_m_axis_tdata[7167:6656]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_13_bits_tkeep = xbar_m_axis_tkeep[847:832]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_13_bits_tlast = xbar_m_axis_tlast[13]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_14_valid = xbar_m_axis_tvalid[14]; // @[BFS.scala 973:40]
  assign io_pe_out_14_bits_tdata = xbar_m_axis_tdata[7679:7168]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_14_bits_tkeep = xbar_m_axis_tkeep[911:896]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_14_bits_tlast = xbar_m_axis_tlast[14]; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_15_valid = xbar_m_axis_tvalid[15]; // @[BFS.scala 973:40]
  assign io_pe_out_15_bits_tdata = xbar_m_axis_tdata[8191:7680]; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_15_bits_tkeep = xbar_m_axis_tkeep[975:960]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_15_bits_tlast = xbar_m_axis_tlast[15]; // @[nf_arm_doce_top.scala 126:21]
  assign xbar_aclk = clock; // @[BFS.scala 968:31]
  assign xbar_aresetn = ~reset; // @[BFS.scala 969:22]
  assign xbar_s_axis_tdata = fat_vertex_filter_io_ddr_out_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign xbar_s_axis_tkeep = {{48'd0}, fat_vertex_filter_io_ddr_out_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign xbar_s_axis_tvalid = fat_vertex_filter_io_ddr_out_valid; // @[BFS.scala 964:27]
  assign xbar_s_axis_tlast = fat_vertex_filter_io_ddr_out_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign xbar_s_axis_tid = 1'h0;
  assign xbar_m_axis_tready = {xbar_io_m_axis_tready_hi,xbar_io_m_axis_tready_lo}; // @[BFS.scala 978:12]
  assign combiner_aclk = clock; // @[BFS.scala 939:37]
  assign combiner_aresetn = ~reset; // @[BFS.scala 940:28]
  assign combiner_s_axis_tdata = {combiner_io_s_axis_tdata_hi,combiner_io_s_axis_tdata_lo}; // @[BFS.scala 941:98]
  assign combiner_s_axis_tkeep = {{48'd0}, _combiner_io_s_axis_tkeep_T_32}; // @[BFS.scala 943:35]
  assign combiner_s_axis_tvalid = {combiner_io_s_axis_tvalid_lo,combiner_io_s_axis_tvalid_lo}; // @[BFS.scala 945:111]
  assign combiner_s_axis_tlast = {combiner_io_s_axis_tlast_hi,combiner_io_s_axis_tlast_lo}; // @[BFS.scala 944:98]
  assign combiner_s_axis_tid = 4'h0;
  assign combiner_m_axis_tready = buffer0_s_axis_tready; // @[BFS.scala 953:23]
  assign buffer0_s_axis_aclk = clock; // @[BFS.scala 951:43]
  assign buffer0_s_axis_aresetn = ~reset; // @[BFS.scala 952:34]
  assign buffer0_s_axis_tdata = combiner_m_axis_tdata; // @[BFS.scala 953:23]
  assign buffer0_s_axis_tkeep = combiner_m_axis_tkeep; // @[BFS.scala 953:23]
  assign buffer0_s_axis_tvalid = combiner_m_axis_tvalid; // @[BFS.scala 953:23]
  assign buffer0_s_axis_tlast = combiner_m_axis_tlast; // @[BFS.scala 953:23]
  assign buffer0_s_axis_tid = combiner_m_axis_tid; // @[BFS.scala 953:23]
  assign buffer0_m_axis_tready = fat_vertex_filter_io_xbar_in_ready; // @[BFS.scala 961:30]
  assign fat_vertex_filter_clock = clock;
  assign fat_vertex_filter_reset = reset;
  assign fat_vertex_filter_io_xbar_in_valid = buffer0_m_axis_tvalid; // @[BFS.scala 959:40]
  assign fat_vertex_filter_io_xbar_in_bits_tdata = buffer0_m_axis_tdata; // @[BFS.scala 956:45]
  assign fat_vertex_filter_io_xbar_in_bits_tkeep = _fat_vertex_filter_io_xbar_in_bits_tkeep_T_128[15:0]; // @[BFS.scala 957:45]
  assign fat_vertex_filter_io_xbar_in_bits_tlast = buffer0_m_axis_tlast; // @[BFS.scala 960:45]
  assign fat_vertex_filter_io_ddr_out_ready = xbar_s_axis_tready; // @[BFS.scala 965:40]
endmodule
module BFS_ps(
  input          clock,
  input          reset,
  input  [63:0]  io_config_awaddr,
  input          io_config_awvalid,
  output         io_config_awready,
  input  [63:0]  io_config_araddr,
  input          io_config_arvalid,
  output         io_config_arready,
  input  [31:0]  io_config_wdata,
  input  [3:0]   io_config_wstrb,
  input          io_config_wvalid,
  output         io_config_wready,
  output [31:0]  io_config_rdata,
  output [1:0]   io_config_rresp,
  output         io_config_rvalid,
  input          io_config_rready,
  output [1:0]   io_config_bresp,
  output         io_config_bvalid,
  input          io_config_bready,
  input          io_PLmemory_0_aw_ready,
  output         io_PLmemory_0_aw_valid,
  output [63:0]  io_PLmemory_0_aw_bits_awaddr,
  output [6:0]   io_PLmemory_0_aw_bits_awid,
  output [7:0]   io_PLmemory_0_aw_bits_awlen,
  output [2:0]   io_PLmemory_0_aw_bits_awsize,
  output [1:0]   io_PLmemory_0_aw_bits_awburst,
  output         io_PLmemory_0_aw_bits_awlock,
  input          io_PLmemory_0_ar_ready,
  output         io_PLmemory_0_ar_valid,
  output [63:0]  io_PLmemory_0_ar_bits_araddr,
  output [6:0]   io_PLmemory_0_ar_bits_arid,
  output [7:0]   io_PLmemory_0_ar_bits_arlen,
  output [2:0]   io_PLmemory_0_ar_bits_arsize,
  output [1:0]   io_PLmemory_0_ar_bits_arburst,
  output         io_PLmemory_0_ar_bits_arlock,
  input          io_PLmemory_0_w_ready,
  output         io_PLmemory_0_w_valid,
  output [511:0] io_PLmemory_0_w_bits_wdata,
  output [63:0]  io_PLmemory_0_w_bits_wstrb,
  output         io_PLmemory_0_w_bits_wlast,
  output         io_PLmemory_0_r_ready,
  input          io_PLmemory_0_r_valid,
  input  [511:0] io_PLmemory_0_r_bits_rdata,
  input  [6:0]   io_PLmemory_0_r_bits_rid,
  input          io_PLmemory_0_r_bits_rlast,
  output         io_PLmemory_0_b_ready,
  input          io_PLmemory_0_b_valid,
  input  [1:0]   io_PLmemory_0_b_bits_bresp,
  input  [6:0]   io_PLmemory_0_b_bits_bid,
  input          io_PLmemory_1_aw_ready,
  output         io_PLmemory_1_aw_valid,
  output [63:0]  io_PLmemory_1_aw_bits_awaddr,
  output [6:0]   io_PLmemory_1_aw_bits_awid,
  output [7:0]   io_PLmemory_1_aw_bits_awlen,
  output [2:0]   io_PLmemory_1_aw_bits_awsize,
  output [1:0]   io_PLmemory_1_aw_bits_awburst,
  output         io_PLmemory_1_aw_bits_awlock,
  input          io_PLmemory_1_ar_ready,
  output         io_PLmemory_1_ar_valid,
  output [63:0]  io_PLmemory_1_ar_bits_araddr,
  output [6:0]   io_PLmemory_1_ar_bits_arid,
  output [7:0]   io_PLmemory_1_ar_bits_arlen,
  output [2:0]   io_PLmemory_1_ar_bits_arsize,
  output [1:0]   io_PLmemory_1_ar_bits_arburst,
  output         io_PLmemory_1_ar_bits_arlock,
  input          io_PLmemory_1_w_ready,
  output         io_PLmemory_1_w_valid,
  output [511:0] io_PLmemory_1_w_bits_wdata,
  output [63:0]  io_PLmemory_1_w_bits_wstrb,
  output         io_PLmemory_1_w_bits_wlast,
  output         io_PLmemory_1_r_ready,
  input          io_PLmemory_1_r_valid,
  input  [511:0] io_PLmemory_1_r_bits_rdata,
  input  [6:0]   io_PLmemory_1_r_bits_rid,
  input          io_PLmemory_1_r_bits_rlast,
  output         io_PLmemory_1_b_ready,
  input          io_PLmemory_1_b_valid,
  input  [1:0]   io_PLmemory_1_b_bits_bresp,
  input  [6:0]   io_PLmemory_1_b_bits_bid,
  input          io_PSmemory_0_aw_ready,
  output         io_PSmemory_0_aw_valid,
  output [63:0]  io_PSmemory_0_aw_bits_awaddr,
  output [5:0]   io_PSmemory_0_aw_bits_awid,
  output [7:0]   io_PSmemory_0_aw_bits_awlen,
  output [2:0]   io_PSmemory_0_aw_bits_awsize,
  output [1:0]   io_PSmemory_0_aw_bits_awburst,
  output         io_PSmemory_0_aw_bits_awlock,
  input          io_PSmemory_0_ar_ready,
  output         io_PSmemory_0_ar_valid,
  output [63:0]  io_PSmemory_0_ar_bits_araddr,
  output [5:0]   io_PSmemory_0_ar_bits_arid,
  output [7:0]   io_PSmemory_0_ar_bits_arlen,
  output [2:0]   io_PSmemory_0_ar_bits_arsize,
  output [1:0]   io_PSmemory_0_ar_bits_arburst,
  output         io_PSmemory_0_ar_bits_arlock,
  input          io_PSmemory_0_w_ready,
  output         io_PSmemory_0_w_valid,
  output [127:0] io_PSmemory_0_w_bits_wdata,
  output [15:0]  io_PSmemory_0_w_bits_wstrb,
  output         io_PSmemory_0_w_bits_wlast,
  output         io_PSmemory_0_r_ready,
  input          io_PSmemory_0_r_valid,
  input  [127:0] io_PSmemory_0_r_bits_rdata,
  input  [5:0]   io_PSmemory_0_r_bits_rid,
  input          io_PSmemory_0_r_bits_rlast,
  output         io_PSmemory_0_b_ready,
  input          io_PSmemory_0_b_valid,
  input  [1:0]   io_PSmemory_0_b_bits_bresp,
  input  [5:0]   io_PSmemory_0_b_bits_bid,
  input          io_PSmemory_1_aw_ready,
  output         io_PSmemory_1_aw_valid,
  output [63:0]  io_PSmemory_1_aw_bits_awaddr,
  output [5:0]   io_PSmemory_1_aw_bits_awid,
  output [7:0]   io_PSmemory_1_aw_bits_awlen,
  output [2:0]   io_PSmemory_1_aw_bits_awsize,
  output [1:0]   io_PSmemory_1_aw_bits_awburst,
  output         io_PSmemory_1_aw_bits_awlock,
  input          io_PSmemory_1_ar_ready,
  output         io_PSmemory_1_ar_valid,
  output [63:0]  io_PSmemory_1_ar_bits_araddr,
  output [5:0]   io_PSmemory_1_ar_bits_arid,
  output [7:0]   io_PSmemory_1_ar_bits_arlen,
  output [2:0]   io_PSmemory_1_ar_bits_arsize,
  output [1:0]   io_PSmemory_1_ar_bits_arburst,
  output         io_PSmemory_1_ar_bits_arlock,
  input          io_PSmemory_1_w_ready,
  output         io_PSmemory_1_w_valid,
  output [127:0] io_PSmemory_1_w_bits_wdata,
  output [15:0]  io_PSmemory_1_w_bits_wstrb,
  output         io_PSmemory_1_w_bits_wlast,
  output         io_PSmemory_1_r_ready,
  input          io_PSmemory_1_r_valid,
  input  [127:0] io_PSmemory_1_r_bits_rdata,
  input  [5:0]   io_PSmemory_1_r_bits_rid,
  input          io_PSmemory_1_r_bits_rlast,
  output         io_PSmemory_1_b_ready,
  input          io_PSmemory_1_b_valid,
  input  [1:0]   io_PSmemory_1_b_bits_bresp,
  input  [5:0]   io_PSmemory_1_b_bits_bid,
  input          io_PSmemory_2_aw_ready,
  output         io_PSmemory_2_aw_valid,
  output [63:0]  io_PSmemory_2_aw_bits_awaddr,
  output [5:0]   io_PSmemory_2_aw_bits_awid,
  output [7:0]   io_PSmemory_2_aw_bits_awlen,
  output [2:0]   io_PSmemory_2_aw_bits_awsize,
  output [1:0]   io_PSmemory_2_aw_bits_awburst,
  output         io_PSmemory_2_aw_bits_awlock,
  input          io_PSmemory_2_ar_ready,
  output         io_PSmemory_2_ar_valid,
  output [63:0]  io_PSmemory_2_ar_bits_araddr,
  output [5:0]   io_PSmemory_2_ar_bits_arid,
  output [7:0]   io_PSmemory_2_ar_bits_arlen,
  output [2:0]   io_PSmemory_2_ar_bits_arsize,
  output [1:0]   io_PSmemory_2_ar_bits_arburst,
  output         io_PSmemory_2_ar_bits_arlock,
  input          io_PSmemory_2_w_ready,
  output         io_PSmemory_2_w_valid,
  output [127:0] io_PSmemory_2_w_bits_wdata,
  output [15:0]  io_PSmemory_2_w_bits_wstrb,
  output         io_PSmemory_2_w_bits_wlast,
  output         io_PSmemory_2_r_ready,
  input          io_PSmemory_2_r_valid,
  input  [127:0] io_PSmemory_2_r_bits_rdata,
  input  [5:0]   io_PSmemory_2_r_bits_rid,
  input          io_PSmemory_2_r_bits_rlast,
  output         io_PSmemory_2_b_ready,
  input          io_PSmemory_2_b_valid,
  input  [1:0]   io_PSmemory_2_b_bits_bresp,
  input  [5:0]   io_PSmemory_2_b_bits_bid,
  input          io_PSmemory_3_aw_ready,
  output         io_PSmemory_3_aw_valid,
  output [63:0]  io_PSmemory_3_aw_bits_awaddr,
  output [5:0]   io_PSmemory_3_aw_bits_awid,
  output [7:0]   io_PSmemory_3_aw_bits_awlen,
  output [2:0]   io_PSmemory_3_aw_bits_awsize,
  output [1:0]   io_PSmemory_3_aw_bits_awburst,
  output         io_PSmemory_3_aw_bits_awlock,
  input          io_PSmemory_3_ar_ready,
  output         io_PSmemory_3_ar_valid,
  output [63:0]  io_PSmemory_3_ar_bits_araddr,
  output [5:0]   io_PSmemory_3_ar_bits_arid,
  output [7:0]   io_PSmemory_3_ar_bits_arlen,
  output [2:0]   io_PSmemory_3_ar_bits_arsize,
  output [1:0]   io_PSmemory_3_ar_bits_arburst,
  output         io_PSmemory_3_ar_bits_arlock,
  input          io_PSmemory_3_w_ready,
  output         io_PSmemory_3_w_valid,
  output [127:0] io_PSmemory_3_w_bits_wdata,
  output [15:0]  io_PSmemory_3_w_bits_wstrb,
  output         io_PSmemory_3_w_bits_wlast,
  output         io_PSmemory_3_r_ready,
  input          io_PSmemory_3_r_valid,
  input  [127:0] io_PSmemory_3_r_bits_rdata,
  input  [5:0]   io_PSmemory_3_r_bits_rid,
  input          io_PSmemory_3_r_bits_rlast,
  output         io_PSmemory_3_b_ready,
  input          io_PSmemory_3_b_valid,
  input  [1:0]   io_PSmemory_3_b_bits_bresp,
  input  [5:0]   io_PSmemory_3_b_bits_bid,
  input          io_Re_memory_out_aw_ready,
  output         io_Re_memory_out_aw_valid,
  output [63:0]  io_Re_memory_out_aw_bits_awaddr,
  output [5:0]   io_Re_memory_out_aw_bits_awid,
  output [7:0]   io_Re_memory_out_aw_bits_awlen,
  output [2:0]   io_Re_memory_out_aw_bits_awsize,
  output [1:0]   io_Re_memory_out_aw_bits_awburst,
  output         io_Re_memory_out_aw_bits_awlock,
  input          io_Re_memory_out_ar_ready,
  output         io_Re_memory_out_ar_valid,
  output [63:0]  io_Re_memory_out_ar_bits_araddr,
  output [5:0]   io_Re_memory_out_ar_bits_arid,
  output [7:0]   io_Re_memory_out_ar_bits_arlen,
  output [2:0]   io_Re_memory_out_ar_bits_arsize,
  output [1:0]   io_Re_memory_out_ar_bits_arburst,
  output         io_Re_memory_out_ar_bits_arlock,
  input          io_Re_memory_out_w_ready,
  output         io_Re_memory_out_w_valid,
  output [511:0] io_Re_memory_out_w_bits_wdata,
  output [63:0]  io_Re_memory_out_w_bits_wstrb,
  output         io_Re_memory_out_w_bits_wlast,
  output         io_Re_memory_out_r_ready,
  input          io_Re_memory_out_r_valid,
  input  [511:0] io_Re_memory_out_r_bits_rdata,
  input  [5:0]   io_Re_memory_out_r_bits_rid,
  input          io_Re_memory_out_r_bits_rlast,
  output         io_Re_memory_out_b_ready,
  input          io_Re_memory_out_b_valid,
  input  [1:0]   io_Re_memory_out_b_bits_bresp,
  input  [5:0]   io_Re_memory_out_b_bits_bid,
  output         io_Re_memory_in_aw_ready,
  input          io_Re_memory_in_aw_valid,
  input  [63:0]  io_Re_memory_in_aw_bits_awaddr,
  input  [9:0]   io_Re_memory_in_aw_bits_awid,
  input  [7:0]   io_Re_memory_in_aw_bits_awlen,
  input  [2:0]   io_Re_memory_in_aw_bits_awsize,
  input  [1:0]   io_Re_memory_in_aw_bits_awburst,
  input          io_Re_memory_in_aw_bits_awlock,
  output         io_Re_memory_in_ar_ready,
  input          io_Re_memory_in_ar_valid,
  input  [63:0]  io_Re_memory_in_ar_bits_araddr,
  input  [9:0]   io_Re_memory_in_ar_bits_arid,
  input  [7:0]   io_Re_memory_in_ar_bits_arlen,
  input  [2:0]   io_Re_memory_in_ar_bits_arsize,
  input  [1:0]   io_Re_memory_in_ar_bits_arburst,
  input          io_Re_memory_in_ar_bits_arlock,
  output         io_Re_memory_in_w_ready,
  input          io_Re_memory_in_w_valid,
  input  [511:0] io_Re_memory_in_w_bits_wdata,
  input  [63:0]  io_Re_memory_in_w_bits_wstrb,
  input          io_Re_memory_in_w_bits_wlast,
  input          io_Re_memory_in_r_ready,
  output         io_Re_memory_in_r_valid,
  output [511:0] io_Re_memory_in_r_bits_rdata,
  output [9:0]   io_Re_memory_in_r_bits_rid,
  output         io_Re_memory_in_r_bits_rlast,
  input          io_Re_memory_in_b_ready,
  output         io_Re_memory_in_b_valid,
  output [1:0]   io_Re_memory_in_b_bits_bresp,
  output [9:0]   io_Re_memory_in_b_bits_bid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  controls_clock; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_reset; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_0; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_1; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_2; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_3; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_4; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_5; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_6; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_7; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_8; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_9; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_10; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_11; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_0; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_1; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_2; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_3; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_4; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_5; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_6; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_7; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_8; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_9; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_10; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_11; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_12; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_13; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_14; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_15; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_signal; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_start; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_level; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_unvisited_size; // @[nf_arm_doce_top_main.scala 30:24]
  wire [63:0] controls_io_traveled_edges; // @[nf_arm_doce_top_main.scala 30:24]
  wire [63:0] controls_io_config_awaddr; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_awvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_awready; // @[nf_arm_doce_top_main.scala 30:24]
  wire [63:0] controls_io_config_araddr; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_arvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_arready; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_config_wdata; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_wvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_wready; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_config_rdata; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_rvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_rready; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_bvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_bready; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_flush_cache; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_flush_cache_end; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 30:24]
  wire  MemController_clock; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_reset; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_out_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_out_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [511:0] MemController_io_cacheable_out_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire [15:0] MemController_io_cacheable_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_0_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_0_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_0_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_1_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_1_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_1_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_2_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_2_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_2_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_3_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_3_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_3_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_4_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_4_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_4_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_5_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_5_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_5_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_6_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_6_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_6_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_7_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_7_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_7_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_8_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_8_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_8_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_9_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_9_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_9_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_10_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_10_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_10_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_11_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_11_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_11_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_12_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_12_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_12_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_13_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_13_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_13_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_14_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_14_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_14_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_15_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_cacheable_in_15_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_cacheable_in_15_bits_tdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_ddr_out_0_aw_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_ddr_out_0_aw_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [63:0] MemController_io_ddr_out_0_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_ddr_out_0_ar_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_ddr_out_0_ar_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [63:0] MemController_io_ddr_out_0_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_ddr_out_0_w_ready; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_ddr_out_0_w_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [511:0] MemController_io_ddr_out_0_w_bits_wdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_ddr_out_0_w_bits_wlast; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_ddr_out_0_r_valid; // @[nf_arm_doce_top_main.scala 33:29]
  wire [511:0] MemController_io_ddr_out_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_ddr_out_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 33:29]
  wire [63:0] MemController_io_tiers_base_addr_0; // @[nf_arm_doce_top_main.scala 33:29]
  wire [63:0] MemController_io_tiers_base_addr_1; // @[nf_arm_doce_top_main.scala 33:29]
  wire [31:0] MemController_io_unvisited_size; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_start; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_signal; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_end; // @[nf_arm_doce_top_main.scala 33:29]
  wire  MemController_io_signal_ack; // @[nf_arm_doce_top_main.scala 33:29]
  wire  Applys_0_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_0_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_0_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_0_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_0_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_0_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_0_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_0_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_0_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_0_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_1_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_1_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_1_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_1_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_1_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_1_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_1_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_1_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_1_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_1_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_2_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_2_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_2_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_2_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_2_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_2_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_2_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_2_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_2_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_2_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_3_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_3_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_3_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_3_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_3_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_3_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_3_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_3_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_3_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_3_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_4_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_4_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_4_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_4_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_4_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_4_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_4_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_4_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_4_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_4_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_4_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_5_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_5_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_5_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_5_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_5_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_5_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_5_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_5_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_5_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_5_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_5_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_6_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_6_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_6_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_6_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_6_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_6_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_6_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_6_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_6_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_6_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_6_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_7_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_7_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_7_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_7_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_7_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_7_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_7_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_7_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_7_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_7_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_7_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_8_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_8_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_8_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_8_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_8_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_8_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_8_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_8_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_8_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_8_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_8_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_9_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_9_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_9_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_9_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_9_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_9_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_9_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_9_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_9_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_9_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_9_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_10_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_10_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_10_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_10_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_10_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_10_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_10_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_10_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_10_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_10_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_10_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_11_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_11_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_11_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_11_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_11_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_11_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_11_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_11_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_11_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_11_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_11_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_12_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_12_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_12_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_12_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_12_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_12_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_12_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_12_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_12_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_12_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_12_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_13_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_13_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_13_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_13_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_13_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_13_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_13_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_13_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_13_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_13_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_13_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_14_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_14_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_14_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_14_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_14_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_14_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_14_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_14_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_14_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_14_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_14_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_15_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_15_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_15_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_15_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Applys_15_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Applys_15_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_15_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_15_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_15_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Applys_15_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Applys_15_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Gathers_clock; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_reset; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_ddr_in_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_ddr_in_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [511:0] Gathers_io_ddr_in_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire [15:0] Gathers_io_ddr_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_0_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_0_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [31:0] Gathers_io_gather_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_1_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_1_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [31:0] Gathers_io_gather_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_2_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_2_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [31:0] Gathers_io_gather_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_3_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_3_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [31:0] Gathers_io_gather_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_level_cache_out_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_level_cache_out_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [511:0] Gathers_io_level_cache_out_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire [15:0] Gathers_io_level_cache_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_level_cache_out_bits_tlast; // @[nf_arm_doce_top_main.scala 37:23]
  wire  LevelCache_clock; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_reset; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_0_ddr_aw_ready; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_0_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 38:26]
  wire [63:0] LevelCache_io_axi_0_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 38:26]
  wire [5:0] LevelCache_io_axi_0_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_0_ddr_w_ready; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_0_ddr_w_valid; // @[nf_arm_doce_top_main.scala 38:26]
  wire [127:0] LevelCache_io_axi_0_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 38:26]
  wire [15:0] LevelCache_io_axi_0_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_1_ddr_aw_ready; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_1_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 38:26]
  wire [63:0] LevelCache_io_axi_1_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 38:26]
  wire [5:0] LevelCache_io_axi_1_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_1_ddr_w_ready; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_1_ddr_w_valid; // @[nf_arm_doce_top_main.scala 38:26]
  wire [127:0] LevelCache_io_axi_1_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 38:26]
  wire [15:0] LevelCache_io_axi_1_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_2_ddr_aw_ready; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_2_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 38:26]
  wire [63:0] LevelCache_io_axi_2_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 38:26]
  wire [5:0] LevelCache_io_axi_2_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_2_ddr_w_ready; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_2_ddr_w_valid; // @[nf_arm_doce_top_main.scala 38:26]
  wire [127:0] LevelCache_io_axi_2_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 38:26]
  wire [15:0] LevelCache_io_axi_2_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_3_ddr_aw_ready; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_3_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 38:26]
  wire [63:0] LevelCache_io_axi_3_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 38:26]
  wire [5:0] LevelCache_io_axi_3_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_3_ddr_w_ready; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_axi_3_ddr_w_valid; // @[nf_arm_doce_top_main.scala 38:26]
  wire [127:0] LevelCache_io_axi_3_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 38:26]
  wire [15:0] LevelCache_io_axi_3_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 38:26]
  wire [511:0] LevelCache_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 38:26]
  wire [63:0] LevelCache_io_gather_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_gather_in_bits_tlast; // @[nf_arm_doce_top_main.scala 38:26]
  wire [31:0] LevelCache_io_level; // @[nf_arm_doce_top_main.scala 38:26]
  wire [63:0] LevelCache_io_level_base_addr; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_end; // @[nf_arm_doce_top_main.scala 38:26]
  wire  LevelCache_io_flush; // @[nf_arm_doce_top_main.scala 38:26]
  wire  Scatters_0_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_0_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Scatters_0_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [7:0] Scatters_0_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 40:16]
  wire [2:0] Scatters_0_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Scatters_0_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Scatters_0_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Scatters_0_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Scatters_0_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Scatters_0_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_0_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_0_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_signal; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_0_io_traveled_edges; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_start; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Scatters_0_io_root; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_0_io_issue_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Scatters_0_io_recv_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_1_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Scatters_1_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [7:0] Scatters_1_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 40:16]
  wire [2:0] Scatters_1_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Scatters_1_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Scatters_1_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Scatters_1_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Scatters_1_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Scatters_1_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_1_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_1_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_signal; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_1_io_traveled_edges; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_1_io_issue_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Scatters_1_io_recv_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_2_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Scatters_2_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [7:0] Scatters_2_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 40:16]
  wire [2:0] Scatters_2_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Scatters_2_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Scatters_2_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Scatters_2_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Scatters_2_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Scatters_2_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_2_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_2_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_signal; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_2_io_traveled_edges; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_2_io_issue_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Scatters_2_io_recv_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_3_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Scatters_3_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [7:0] Scatters_3_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 40:16]
  wire [2:0] Scatters_3_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Scatters_3_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Scatters_3_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Scatters_3_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Scatters_3_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Scatters_3_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_3_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_3_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_signal; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Scatters_3_io_traveled_edges; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Scatters_3_io_issue_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Scatters_3_io_recv_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcaster_clock; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_reset; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_0_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_0_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [127:0] Broadcaster_io_ddr_in_0_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [3:0] Broadcaster_io_ddr_in_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_0_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_1_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_1_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [127:0] Broadcaster_io_ddr_in_1_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [3:0] Broadcaster_io_ddr_in_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_1_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_2_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_2_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [127:0] Broadcaster_io_ddr_in_2_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [3:0] Broadcaster_io_ddr_in_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_2_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_3_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_3_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [127:0] Broadcaster_io_ddr_in_3_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [3:0] Broadcaster_io_ddr_in_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_ddr_in_3_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_0_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_0_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_0_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_1_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_1_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_1_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_2_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_2_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_2_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_3_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_3_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_3_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_4_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_4_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_4_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_4_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_5_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_5_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_5_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_5_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_5_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_6_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_6_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_6_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_6_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_6_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_7_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_7_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_7_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_7_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_7_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_8_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_8_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_8_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_8_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_8_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_9_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_9_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_9_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_9_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_9_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_10_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_10_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_10_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_10_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_10_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_11_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_11_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_11_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_11_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_11_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_12_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_12_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_12_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_12_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_12_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_13_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_13_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_13_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_13_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_13_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_14_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_14_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_14_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_14_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_14_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_15_ready; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_15_valid; // @[nf_arm_doce_top_main.scala 43:27]
  wire [511:0] Broadcaster_io_pe_out_15_bits_tdata; // @[nf_arm_doce_top_main.scala 43:27]
  wire [15:0] Broadcaster_io_pe_out_15_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:27]
  wire  Broadcaster_io_pe_out_15_bits_tlast; // @[nf_arm_doce_top_main.scala 43:27]
  wire  _T_1 = ~io_PSmemory_0_r_valid; // @[nf_arm_doce_top_main.scala 45:77]
  wire  _T_2 = LevelCache_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 46:35]
  wire  _T_3 = ~io_PSmemory_0_r_valid & _T_2; // @[nf_arm_doce_top_main.scala 45:89]
  wire  _T_5 = _T_3 & ~LevelCache_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 46:46]
    (*dont_touch = "true" *)reg [30:0] ar_ready_counter1; // @[Counter.scala 60:40]
  wire  wrap_wrap = ar_ready_counter1 == 31'h7ffffffe; // @[Counter.scala 72:24]
  wire [30:0] _wrap_value_T_1 = ar_ready_counter1 + 31'h1; // @[Counter.scala 76:24]
    (*dont_touch = "true" *)reg [31:0] axi_ready_counter_0; // @[nf_arm_doce_top_main.scala 49:34]
    (*dont_touch = "true" *)reg [31:0] axi_ready_counter_1; // @[nf_arm_doce_top_main.scala 49:34]
    (*dont_touch = "true" *)reg [31:0] axi_ready_counter_2; // @[nf_arm_doce_top_main.scala 49:34]
    (*dont_touch = "true" *)reg [31:0] axi_ready_counter_3; // @[nf_arm_doce_top_main.scala 49:34]
  wire  _T_9 = ~io_PSmemory_0_ar_valid; // @[nf_arm_doce_top_main.scala 54:32]
  wire  _T_10 = ~io_PSmemory_0_w_valid & _T_1 & _T_9; // @[nf_arm_doce_top_main.scala 53:84]
  wire  _T_12 = _T_10 & ~io_PSmemory_0_aw_valid; // @[nf_arm_doce_top_main.scala 54:44]
  wire  _T_13 = Gathers_io_ddr_in_valid; // @[nf_arm_doce_top_main.scala 55:32]
  wire  _T_14 = _T_10 & ~io_PSmemory_0_aw_valid & _T_13; // @[nf_arm_doce_top_main.scala 54:83]
  wire [31:0] _axi_ready_counter_0_T_1 = axi_ready_counter_0 + 32'h1; // @[nf_arm_doce_top_main.scala 56:15]
  wire  _T_15 = ~io_PSmemory_1_w_valid; // @[nf_arm_doce_top_main.scala 53:34]
  wire  _T_16 = ~io_PSmemory_1_r_valid; // @[nf_arm_doce_top_main.scala 53:72]
  wire  _T_18 = ~io_PSmemory_1_ar_valid; // @[nf_arm_doce_top_main.scala 54:32]
  wire  _T_19 = ~io_PSmemory_1_w_valid & ~io_PSmemory_1_r_valid & _T_18; // @[nf_arm_doce_top_main.scala 53:84]
  wire  _T_20 = ~io_PSmemory_1_aw_valid; // @[nf_arm_doce_top_main.scala 54:71]
  wire  _T_23 = _T_19 & ~io_PSmemory_1_aw_valid & _T_13; // @[nf_arm_doce_top_main.scala 54:83]
  wire [31:0] _axi_ready_counter_1_T_1 = axi_ready_counter_1 + 32'h1; // @[nf_arm_doce_top_main.scala 56:15]
  wire  _T_24 = ~io_PSmemory_2_w_valid; // @[nf_arm_doce_top_main.scala 53:34]
  wire  _T_25 = ~io_PSmemory_2_r_valid; // @[nf_arm_doce_top_main.scala 53:72]
  wire  _T_27 = ~io_PSmemory_2_ar_valid; // @[nf_arm_doce_top_main.scala 54:32]
  wire  _T_28 = ~io_PSmemory_2_w_valid & ~io_PSmemory_2_r_valid & _T_27; // @[nf_arm_doce_top_main.scala 53:84]
  wire  _T_29 = ~io_PSmemory_2_aw_valid; // @[nf_arm_doce_top_main.scala 54:71]
  wire  _T_32 = _T_28 & ~io_PSmemory_2_aw_valid & _T_13; // @[nf_arm_doce_top_main.scala 54:83]
  wire [31:0] _axi_ready_counter_2_T_1 = axi_ready_counter_2 + 32'h1; // @[nf_arm_doce_top_main.scala 56:15]
  wire  _T_33 = ~io_PSmemory_3_w_valid; // @[nf_arm_doce_top_main.scala 53:34]
  wire  _T_34 = ~io_PSmemory_3_r_valid; // @[nf_arm_doce_top_main.scala 53:72]
  wire  _T_36 = ~io_PSmemory_3_ar_valid; // @[nf_arm_doce_top_main.scala 54:32]
  wire  _T_37 = ~io_PSmemory_3_w_valid & ~io_PSmemory_3_r_valid & _T_36; // @[nf_arm_doce_top_main.scala 53:84]
  wire  _T_38 = ~io_PSmemory_3_aw_valid; // @[nf_arm_doce_top_main.scala 54:71]
  wire  _T_41 = _T_37 & ~io_PSmemory_3_aw_valid & _T_13; // @[nf_arm_doce_top_main.scala 54:83]
  wire [31:0] _axi_ready_counter_3_T_1 = axi_ready_counter_3 + 32'h1; // @[nf_arm_doce_top_main.scala 56:15]
    (*dont_touch = "true" *)reg [31:0] axi_all_ready_counter; // @[nf_arm_doce_top_main.scala 60:38]
  wire  _T_50 = _T_12 & _T_15; // @[nf_arm_doce_top_main.scala 63:80]
  wire  _T_54 = _T_50 & _T_16 & _T_18; // @[nf_arm_doce_top_main.scala 64:78]
  wire  _T_58 = _T_54 & _T_20 & _T_24; // @[nf_arm_doce_top_main.scala 65:80]
  wire  _T_62 = _T_58 & _T_25 & _T_27; // @[nf_arm_doce_top_main.scala 66:78]
  wire  _T_66 = _T_62 & _T_29 & _T_33; // @[nf_arm_doce_top_main.scala 67:80]
  wire  _T_70 = _T_66 & _T_34 & _T_36; // @[nf_arm_doce_top_main.scala 68:78]
  wire  _T_74 = _T_70 & _T_38 & _T_13; // @[nf_arm_doce_top_main.scala 69:80]
  wire [31:0] _axi_all_ready_counter_T_1 = axi_all_ready_counter + 32'h1; // @[nf_arm_doce_top_main.scala 71:52]
    (*dont_touch = "true" *)reg [31:0] axi_r_all_ready_counter; // @[nf_arm_doce_top_main.scala 73:40]
  wire  _T_77 = _T_1 & _T_9; // @[nf_arm_doce_top_main.scala 75:43]
  wire  _T_79 = _T_77 & _T_16; // @[nf_arm_doce_top_main.scala 76:41]
  wire  _T_81 = _T_79 & _T_18; // @[nf_arm_doce_top_main.scala 77:40]
  wire  _T_83 = _T_81 & _T_25; // @[nf_arm_doce_top_main.scala 78:41]
  wire  _T_85 = _T_83 & _T_27; // @[nf_arm_doce_top_main.scala 79:41]
  wire  _T_87 = _T_85 & _T_34; // @[nf_arm_doce_top_main.scala 80:41]
  wire  _T_89 = _T_87 & _T_36; // @[nf_arm_doce_top_main.scala 81:40]
  wire  _T_91 = _T_89 & _T_13; // @[nf_arm_doce_top_main.scala 82:41]
  wire [31:0] _axi_r_all_ready_counter_T_1 = axi_r_all_ready_counter + 32'h1; // @[nf_arm_doce_top_main.scala 84:56]
  wire [63:0] _controls_io_traveled_edges_T_1 = Scatters_0_io_traveled_edges + Scatters_1_io_traveled_edges; // @[nf_arm_doce_top_main.scala 142:80]
  wire [63:0] _controls_io_traveled_edges_T_3 = _controls_io_traveled_edges_T_1 + Scatters_2_io_traveled_edges; // @[nf_arm_doce_top_main.scala 142:80]
  wire  _Scatters_0_io_recv_sync_WIRE_1 = Scatters_1_io_issue_sync; // @[nf_arm_doce_top_main.scala 162:32 nf_arm_doce_top_main.scala 162:32]
  wire  _Scatters_0_io_recv_sync_WIRE_0 = Scatters_0_io_issue_sync; // @[nf_arm_doce_top_main.scala 162:32 nf_arm_doce_top_main.scala 162:32]
  wire [1:0] Scatters_0_io_recv_sync_lo = {_Scatters_0_io_recv_sync_WIRE_1,_Scatters_0_io_recv_sync_WIRE_0}; // @[nf_arm_doce_top_main.scala 162:75]
  wire  _Scatters_0_io_recv_sync_WIRE_3 = Scatters_3_io_issue_sync; // @[nf_arm_doce_top_main.scala 162:32 nf_arm_doce_top_main.scala 162:32]
  wire  _Scatters_0_io_recv_sync_WIRE_2 = Scatters_2_io_issue_sync; // @[nf_arm_doce_top_main.scala 162:32 nf_arm_doce_top_main.scala 162:32]
  wire [1:0] Scatters_0_io_recv_sync_hi = {_Scatters_0_io_recv_sync_WIRE_3,_Scatters_0_io_recv_sync_WIRE_2}; // @[nf_arm_doce_top_main.scala 162:75]
  controller controls ( // @[nf_arm_doce_top_main.scala 30:24]
    .clock(controls_clock),
    .reset(controls_reset),
    .io_data_0(controls_io_data_0),
    .io_data_1(controls_io_data_1),
    .io_data_2(controls_io_data_2),
    .io_data_3(controls_io_data_3),
    .io_data_4(controls_io_data_4),
    .io_data_5(controls_io_data_5),
    .io_data_6(controls_io_data_6),
    .io_data_7(controls_io_data_7),
    .io_data_8(controls_io_data_8),
    .io_data_9(controls_io_data_9),
    .io_data_10(controls_io_data_10),
    .io_data_11(controls_io_data_11),
    .io_fin_0(controls_io_fin_0),
    .io_fin_1(controls_io_fin_1),
    .io_fin_2(controls_io_fin_2),
    .io_fin_3(controls_io_fin_3),
    .io_fin_4(controls_io_fin_4),
    .io_fin_5(controls_io_fin_5),
    .io_fin_6(controls_io_fin_6),
    .io_fin_7(controls_io_fin_7),
    .io_fin_8(controls_io_fin_8),
    .io_fin_9(controls_io_fin_9),
    .io_fin_10(controls_io_fin_10),
    .io_fin_11(controls_io_fin_11),
    .io_fin_12(controls_io_fin_12),
    .io_fin_13(controls_io_fin_13),
    .io_fin_14(controls_io_fin_14),
    .io_fin_15(controls_io_fin_15),
    .io_signal(controls_io_signal),
    .io_start(controls_io_start),
    .io_level(controls_io_level),
    .io_unvisited_size(controls_io_unvisited_size),
    .io_traveled_edges(controls_io_traveled_edges),
    .io_config_awaddr(controls_io_config_awaddr),
    .io_config_awvalid(controls_io_config_awvalid),
    .io_config_awready(controls_io_config_awready),
    .io_config_araddr(controls_io_config_araddr),
    .io_config_arvalid(controls_io_config_arvalid),
    .io_config_arready(controls_io_config_arready),
    .io_config_wdata(controls_io_config_wdata),
    .io_config_wvalid(controls_io_config_wvalid),
    .io_config_wready(controls_io_config_wready),
    .io_config_rdata(controls_io_config_rdata),
    .io_config_rvalid(controls_io_config_rvalid),
    .io_config_rready(controls_io_config_rready),
    .io_config_bvalid(controls_io_config_bvalid),
    .io_config_bready(controls_io_config_bready),
    .io_flush_cache(controls_io_flush_cache),
    .io_flush_cache_end(controls_io_flush_cache_end),
    .io_signal_ack(controls_io_signal_ack)
  );
  multi_port_mc MemController ( // @[nf_arm_doce_top_main.scala 33:29]
    .clock(MemController_clock),
    .reset(MemController_reset),
    .io_cacheable_out_ready(MemController_io_cacheable_out_ready),
    .io_cacheable_out_valid(MemController_io_cacheable_out_valid),
    .io_cacheable_out_bits_tdata(MemController_io_cacheable_out_bits_tdata),
    .io_cacheable_out_bits_tkeep(MemController_io_cacheable_out_bits_tkeep),
    .io_cacheable_in_0_ready(MemController_io_cacheable_in_0_ready),
    .io_cacheable_in_0_valid(MemController_io_cacheable_in_0_valid),
    .io_cacheable_in_0_bits_tdata(MemController_io_cacheable_in_0_bits_tdata),
    .io_cacheable_in_1_ready(MemController_io_cacheable_in_1_ready),
    .io_cacheable_in_1_valid(MemController_io_cacheable_in_1_valid),
    .io_cacheable_in_1_bits_tdata(MemController_io_cacheable_in_1_bits_tdata),
    .io_cacheable_in_2_ready(MemController_io_cacheable_in_2_ready),
    .io_cacheable_in_2_valid(MemController_io_cacheable_in_2_valid),
    .io_cacheable_in_2_bits_tdata(MemController_io_cacheable_in_2_bits_tdata),
    .io_cacheable_in_3_ready(MemController_io_cacheable_in_3_ready),
    .io_cacheable_in_3_valid(MemController_io_cacheable_in_3_valid),
    .io_cacheable_in_3_bits_tdata(MemController_io_cacheable_in_3_bits_tdata),
    .io_cacheable_in_4_ready(MemController_io_cacheable_in_4_ready),
    .io_cacheable_in_4_valid(MemController_io_cacheable_in_4_valid),
    .io_cacheable_in_4_bits_tdata(MemController_io_cacheable_in_4_bits_tdata),
    .io_cacheable_in_5_ready(MemController_io_cacheable_in_5_ready),
    .io_cacheable_in_5_valid(MemController_io_cacheable_in_5_valid),
    .io_cacheable_in_5_bits_tdata(MemController_io_cacheable_in_5_bits_tdata),
    .io_cacheable_in_6_ready(MemController_io_cacheable_in_6_ready),
    .io_cacheable_in_6_valid(MemController_io_cacheable_in_6_valid),
    .io_cacheable_in_6_bits_tdata(MemController_io_cacheable_in_6_bits_tdata),
    .io_cacheable_in_7_ready(MemController_io_cacheable_in_7_ready),
    .io_cacheable_in_7_valid(MemController_io_cacheable_in_7_valid),
    .io_cacheable_in_7_bits_tdata(MemController_io_cacheable_in_7_bits_tdata),
    .io_cacheable_in_8_ready(MemController_io_cacheable_in_8_ready),
    .io_cacheable_in_8_valid(MemController_io_cacheable_in_8_valid),
    .io_cacheable_in_8_bits_tdata(MemController_io_cacheable_in_8_bits_tdata),
    .io_cacheable_in_9_ready(MemController_io_cacheable_in_9_ready),
    .io_cacheable_in_9_valid(MemController_io_cacheable_in_9_valid),
    .io_cacheable_in_9_bits_tdata(MemController_io_cacheable_in_9_bits_tdata),
    .io_cacheable_in_10_ready(MemController_io_cacheable_in_10_ready),
    .io_cacheable_in_10_valid(MemController_io_cacheable_in_10_valid),
    .io_cacheable_in_10_bits_tdata(MemController_io_cacheable_in_10_bits_tdata),
    .io_cacheable_in_11_ready(MemController_io_cacheable_in_11_ready),
    .io_cacheable_in_11_valid(MemController_io_cacheable_in_11_valid),
    .io_cacheable_in_11_bits_tdata(MemController_io_cacheable_in_11_bits_tdata),
    .io_cacheable_in_12_ready(MemController_io_cacheable_in_12_ready),
    .io_cacheable_in_12_valid(MemController_io_cacheable_in_12_valid),
    .io_cacheable_in_12_bits_tdata(MemController_io_cacheable_in_12_bits_tdata),
    .io_cacheable_in_13_ready(MemController_io_cacheable_in_13_ready),
    .io_cacheable_in_13_valid(MemController_io_cacheable_in_13_valid),
    .io_cacheable_in_13_bits_tdata(MemController_io_cacheable_in_13_bits_tdata),
    .io_cacheable_in_14_ready(MemController_io_cacheable_in_14_ready),
    .io_cacheable_in_14_valid(MemController_io_cacheable_in_14_valid),
    .io_cacheable_in_14_bits_tdata(MemController_io_cacheable_in_14_bits_tdata),
    .io_cacheable_in_15_ready(MemController_io_cacheable_in_15_ready),
    .io_cacheable_in_15_valid(MemController_io_cacheable_in_15_valid),
    .io_cacheable_in_15_bits_tdata(MemController_io_cacheable_in_15_bits_tdata),
    .io_ddr_out_0_aw_ready(MemController_io_ddr_out_0_aw_ready),
    .io_ddr_out_0_aw_valid(MemController_io_ddr_out_0_aw_valid),
    .io_ddr_out_0_aw_bits_awaddr(MemController_io_ddr_out_0_aw_bits_awaddr),
    .io_ddr_out_0_ar_ready(MemController_io_ddr_out_0_ar_ready),
    .io_ddr_out_0_ar_valid(MemController_io_ddr_out_0_ar_valid),
    .io_ddr_out_0_ar_bits_araddr(MemController_io_ddr_out_0_ar_bits_araddr),
    .io_ddr_out_0_w_ready(MemController_io_ddr_out_0_w_ready),
    .io_ddr_out_0_w_valid(MemController_io_ddr_out_0_w_valid),
    .io_ddr_out_0_w_bits_wdata(MemController_io_ddr_out_0_w_bits_wdata),
    .io_ddr_out_0_w_bits_wlast(MemController_io_ddr_out_0_w_bits_wlast),
    .io_ddr_out_0_r_valid(MemController_io_ddr_out_0_r_valid),
    .io_ddr_out_0_r_bits_rdata(MemController_io_ddr_out_0_r_bits_rdata),
    .io_ddr_out_0_r_bits_rlast(MemController_io_ddr_out_0_r_bits_rlast),
    .io_tiers_base_addr_0(MemController_io_tiers_base_addr_0),
    .io_tiers_base_addr_1(MemController_io_tiers_base_addr_1),
    .io_unvisited_size(MemController_io_unvisited_size),
    .io_start(MemController_io_start),
    .io_signal(MemController_io_signal),
    .io_end(MemController_io_end),
    .io_signal_ack(MemController_io_signal_ack)
  );
  Scatter Applys_0 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_0_clock),
    .reset(Applys_0_reset),
    .io_xbar_in_ready(Applys_0_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_0_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_0_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_0_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_0_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_0_io_ddr_out_bits_tdata),
    .io_end(Applys_0_io_end)
  );
  Scatter_1 Applys_1 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_1_clock),
    .reset(Applys_1_reset),
    .io_xbar_in_ready(Applys_1_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_1_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_1_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_1_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_1_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_1_io_ddr_out_bits_tdata),
    .io_end(Applys_1_io_end)
  );
  Scatter_2 Applys_2 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_2_clock),
    .reset(Applys_2_reset),
    .io_xbar_in_ready(Applys_2_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_2_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_2_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_2_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_2_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_2_io_ddr_out_bits_tdata),
    .io_end(Applys_2_io_end)
  );
  Scatter_3 Applys_3 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_3_clock),
    .reset(Applys_3_reset),
    .io_xbar_in_ready(Applys_3_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_3_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_3_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_3_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_3_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_3_io_ddr_out_bits_tdata),
    .io_end(Applys_3_io_end)
  );
  Scatter_4 Applys_4 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_4_clock),
    .reset(Applys_4_reset),
    .io_xbar_in_ready(Applys_4_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_4_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_4_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_4_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_4_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_4_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_4_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_4_io_ddr_out_bits_tdata),
    .io_end(Applys_4_io_end)
  );
  Scatter_5 Applys_5 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_5_clock),
    .reset(Applys_5_reset),
    .io_xbar_in_ready(Applys_5_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_5_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_5_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_5_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_5_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_5_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_5_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_5_io_ddr_out_bits_tdata),
    .io_end(Applys_5_io_end)
  );
  Scatter_6 Applys_6 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_6_clock),
    .reset(Applys_6_reset),
    .io_xbar_in_ready(Applys_6_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_6_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_6_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_6_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_6_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_6_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_6_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_6_io_ddr_out_bits_tdata),
    .io_end(Applys_6_io_end)
  );
  Scatter_7 Applys_7 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_7_clock),
    .reset(Applys_7_reset),
    .io_xbar_in_ready(Applys_7_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_7_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_7_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_7_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_7_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_7_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_7_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_7_io_ddr_out_bits_tdata),
    .io_end(Applys_7_io_end)
  );
  Scatter_8 Applys_8 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_8_clock),
    .reset(Applys_8_reset),
    .io_xbar_in_ready(Applys_8_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_8_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_8_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_8_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_8_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_8_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_8_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_8_io_ddr_out_bits_tdata),
    .io_end(Applys_8_io_end)
  );
  Scatter_9 Applys_9 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_9_clock),
    .reset(Applys_9_reset),
    .io_xbar_in_ready(Applys_9_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_9_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_9_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_9_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_9_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_9_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_9_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_9_io_ddr_out_bits_tdata),
    .io_end(Applys_9_io_end)
  );
  Scatter_10 Applys_10 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_10_clock),
    .reset(Applys_10_reset),
    .io_xbar_in_ready(Applys_10_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_10_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_10_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_10_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_10_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_10_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_10_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_10_io_ddr_out_bits_tdata),
    .io_end(Applys_10_io_end)
  );
  Scatter_11 Applys_11 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_11_clock),
    .reset(Applys_11_reset),
    .io_xbar_in_ready(Applys_11_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_11_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_11_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_11_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_11_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_11_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_11_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_11_io_ddr_out_bits_tdata),
    .io_end(Applys_11_io_end)
  );
  Scatter_12 Applys_12 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_12_clock),
    .reset(Applys_12_reset),
    .io_xbar_in_ready(Applys_12_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_12_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_12_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_12_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_12_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_12_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_12_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_12_io_ddr_out_bits_tdata),
    .io_end(Applys_12_io_end)
  );
  Scatter_13 Applys_13 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_13_clock),
    .reset(Applys_13_reset),
    .io_xbar_in_ready(Applys_13_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_13_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_13_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_13_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_13_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_13_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_13_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_13_io_ddr_out_bits_tdata),
    .io_end(Applys_13_io_end)
  );
  Scatter_14 Applys_14 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_14_clock),
    .reset(Applys_14_reset),
    .io_xbar_in_ready(Applys_14_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_14_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_14_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_14_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_14_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_14_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_14_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_14_io_ddr_out_bits_tdata),
    .io_end(Applys_14_io_end)
  );
  Scatter_15 Applys_15 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Applys_15_clock),
    .reset(Applys_15_reset),
    .io_xbar_in_ready(Applys_15_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_15_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_15_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_15_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_15_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(Applys_15_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_15_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_15_io_ddr_out_bits_tdata),
    .io_end(Applys_15_io_end)
  );
  Gather Gathers ( // @[nf_arm_doce_top_main.scala 37:23]
    .clock(Gathers_clock),
    .reset(Gathers_reset),
    .io_ddr_in_ready(Gathers_io_ddr_in_ready),
    .io_ddr_in_valid(Gathers_io_ddr_in_valid),
    .io_ddr_in_bits_tdata(Gathers_io_ddr_in_bits_tdata),
    .io_ddr_in_bits_tkeep(Gathers_io_ddr_in_bits_tkeep),
    .io_gather_out_0_ready(Gathers_io_gather_out_0_ready),
    .io_gather_out_0_valid(Gathers_io_gather_out_0_valid),
    .io_gather_out_0_bits_tdata(Gathers_io_gather_out_0_bits_tdata),
    .io_gather_out_1_ready(Gathers_io_gather_out_1_ready),
    .io_gather_out_1_valid(Gathers_io_gather_out_1_valid),
    .io_gather_out_1_bits_tdata(Gathers_io_gather_out_1_bits_tdata),
    .io_gather_out_2_ready(Gathers_io_gather_out_2_ready),
    .io_gather_out_2_valid(Gathers_io_gather_out_2_valid),
    .io_gather_out_2_bits_tdata(Gathers_io_gather_out_2_bits_tdata),
    .io_gather_out_3_ready(Gathers_io_gather_out_3_ready),
    .io_gather_out_3_valid(Gathers_io_gather_out_3_valid),
    .io_gather_out_3_bits_tdata(Gathers_io_gather_out_3_bits_tdata),
    .io_level_cache_out_ready(Gathers_io_level_cache_out_ready),
    .io_level_cache_out_valid(Gathers_io_level_cache_out_valid),
    .io_level_cache_out_bits_tdata(Gathers_io_level_cache_out_bits_tdata),
    .io_level_cache_out_bits_tkeep(Gathers_io_level_cache_out_bits_tkeep),
    .io_level_cache_out_bits_tlast(Gathers_io_level_cache_out_bits_tlast)
  );
  Apply LevelCache ( // @[nf_arm_doce_top_main.scala 38:26]
    .clock(LevelCache_clock),
    .reset(LevelCache_reset),
    .io_axi_0_ddr_aw_ready(LevelCache_io_axi_0_ddr_aw_ready),
    .io_axi_0_ddr_aw_valid(LevelCache_io_axi_0_ddr_aw_valid),
    .io_axi_0_ddr_aw_bits_awaddr(LevelCache_io_axi_0_ddr_aw_bits_awaddr),
    .io_axi_0_ddr_aw_bits_awid(LevelCache_io_axi_0_ddr_aw_bits_awid),
    .io_axi_0_ddr_w_ready(LevelCache_io_axi_0_ddr_w_ready),
    .io_axi_0_ddr_w_valid(LevelCache_io_axi_0_ddr_w_valid),
    .io_axi_0_ddr_w_bits_wdata(LevelCache_io_axi_0_ddr_w_bits_wdata),
    .io_axi_0_ddr_w_bits_wstrb(LevelCache_io_axi_0_ddr_w_bits_wstrb),
    .io_axi_1_ddr_aw_ready(LevelCache_io_axi_1_ddr_aw_ready),
    .io_axi_1_ddr_aw_valid(LevelCache_io_axi_1_ddr_aw_valid),
    .io_axi_1_ddr_aw_bits_awaddr(LevelCache_io_axi_1_ddr_aw_bits_awaddr),
    .io_axi_1_ddr_aw_bits_awid(LevelCache_io_axi_1_ddr_aw_bits_awid),
    .io_axi_1_ddr_w_ready(LevelCache_io_axi_1_ddr_w_ready),
    .io_axi_1_ddr_w_valid(LevelCache_io_axi_1_ddr_w_valid),
    .io_axi_1_ddr_w_bits_wdata(LevelCache_io_axi_1_ddr_w_bits_wdata),
    .io_axi_1_ddr_w_bits_wstrb(LevelCache_io_axi_1_ddr_w_bits_wstrb),
    .io_axi_2_ddr_aw_ready(LevelCache_io_axi_2_ddr_aw_ready),
    .io_axi_2_ddr_aw_valid(LevelCache_io_axi_2_ddr_aw_valid),
    .io_axi_2_ddr_aw_bits_awaddr(LevelCache_io_axi_2_ddr_aw_bits_awaddr),
    .io_axi_2_ddr_aw_bits_awid(LevelCache_io_axi_2_ddr_aw_bits_awid),
    .io_axi_2_ddr_w_ready(LevelCache_io_axi_2_ddr_w_ready),
    .io_axi_2_ddr_w_valid(LevelCache_io_axi_2_ddr_w_valid),
    .io_axi_2_ddr_w_bits_wdata(LevelCache_io_axi_2_ddr_w_bits_wdata),
    .io_axi_2_ddr_w_bits_wstrb(LevelCache_io_axi_2_ddr_w_bits_wstrb),
    .io_axi_3_ddr_aw_ready(LevelCache_io_axi_3_ddr_aw_ready),
    .io_axi_3_ddr_aw_valid(LevelCache_io_axi_3_ddr_aw_valid),
    .io_axi_3_ddr_aw_bits_awaddr(LevelCache_io_axi_3_ddr_aw_bits_awaddr),
    .io_axi_3_ddr_aw_bits_awid(LevelCache_io_axi_3_ddr_aw_bits_awid),
    .io_axi_3_ddr_w_ready(LevelCache_io_axi_3_ddr_w_ready),
    .io_axi_3_ddr_w_valid(LevelCache_io_axi_3_ddr_w_valid),
    .io_axi_3_ddr_w_bits_wdata(LevelCache_io_axi_3_ddr_w_bits_wdata),
    .io_axi_3_ddr_w_bits_wstrb(LevelCache_io_axi_3_ddr_w_bits_wstrb),
    .io_gather_in_ready(LevelCache_io_gather_in_ready),
    .io_gather_in_valid(LevelCache_io_gather_in_valid),
    .io_gather_in_bits_tdata(LevelCache_io_gather_in_bits_tdata),
    .io_gather_in_bits_tkeep(LevelCache_io_gather_in_bits_tkeep),
    .io_gather_in_bits_tlast(LevelCache_io_gather_in_bits_tlast),
    .io_level(LevelCache_io_level),
    .io_level_base_addr(LevelCache_io_level_base_addr),
    .io_end(LevelCache_io_end),
    .io_flush(LevelCache_io_flush)
  );
  Broadcast Scatters_0 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Scatters_0_clock),
    .reset(Scatters_0_reset),
    .io_ddr_ar_ready(Scatters_0_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_0_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_0_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_0_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_0_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_0_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_0_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_0_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_0_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_0_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_0_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_0_io_gather_in_ready),
    .io_gather_in_valid(Scatters_0_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_0_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_0_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_0_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_0_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_0_io_xbar_out_bits_tkeep),
    .io_xbar_out_bits_tlast(Scatters_0_io_xbar_out_bits_tlast),
    .io_embedding_base_addr(Scatters_0_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_0_io_edge_base_addr),
    .io_signal(Scatters_0_io_signal),
    .io_traveled_edges(Scatters_0_io_traveled_edges),
    .io_start(Scatters_0_io_start),
    .io_root(Scatters_0_io_root),
    .io_issue_sync(Scatters_0_io_issue_sync),
    .io_recv_sync(Scatters_0_io_recv_sync)
  );
  Broadcast_1 Scatters_1 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Scatters_1_clock),
    .reset(Scatters_1_reset),
    .io_ddr_ar_ready(Scatters_1_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_1_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_1_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_1_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_1_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_1_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_1_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_1_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_1_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_1_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_1_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_1_io_gather_in_ready),
    .io_gather_in_valid(Scatters_1_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_1_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_1_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_1_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_1_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_1_io_xbar_out_bits_tkeep),
    .io_xbar_out_bits_tlast(Scatters_1_io_xbar_out_bits_tlast),
    .io_embedding_base_addr(Scatters_1_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_1_io_edge_base_addr),
    .io_signal(Scatters_1_io_signal),
    .io_traveled_edges(Scatters_1_io_traveled_edges),
    .io_issue_sync(Scatters_1_io_issue_sync),
    .io_recv_sync(Scatters_1_io_recv_sync)
  );
  Broadcast_2 Scatters_2 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Scatters_2_clock),
    .reset(Scatters_2_reset),
    .io_ddr_ar_ready(Scatters_2_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_2_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_2_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_2_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_2_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_2_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_2_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_2_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_2_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_2_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_2_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_2_io_gather_in_ready),
    .io_gather_in_valid(Scatters_2_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_2_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_2_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_2_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_2_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_2_io_xbar_out_bits_tkeep),
    .io_xbar_out_bits_tlast(Scatters_2_io_xbar_out_bits_tlast),
    .io_embedding_base_addr(Scatters_2_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_2_io_edge_base_addr),
    .io_signal(Scatters_2_io_signal),
    .io_traveled_edges(Scatters_2_io_traveled_edges),
    .io_issue_sync(Scatters_2_io_issue_sync),
    .io_recv_sync(Scatters_2_io_recv_sync)
  );
  Broadcast_3 Scatters_3 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Scatters_3_clock),
    .reset(Scatters_3_reset),
    .io_ddr_ar_ready(Scatters_3_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_3_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_3_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_3_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_3_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_3_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_3_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_3_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_3_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_3_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_3_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_3_io_gather_in_ready),
    .io_gather_in_valid(Scatters_3_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_3_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_3_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_3_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_3_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_3_io_xbar_out_bits_tkeep),
    .io_xbar_out_bits_tlast(Scatters_3_io_xbar_out_bits_tlast),
    .io_embedding_base_addr(Scatters_3_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_3_io_edge_base_addr),
    .io_signal(Scatters_3_io_signal),
    .io_traveled_edges(Scatters_3_io_traveled_edges),
    .io_issue_sync(Scatters_3_io_issue_sync),
    .io_recv_sync(Scatters_3_io_recv_sync)
  );
  broadcast_xbar Broadcaster ( // @[nf_arm_doce_top_main.scala 43:27]
    .clock(Broadcaster_clock),
    .reset(Broadcaster_reset),
    .io_ddr_in_0_ready(Broadcaster_io_ddr_in_0_ready),
    .io_ddr_in_0_valid(Broadcaster_io_ddr_in_0_valid),
    .io_ddr_in_0_bits_tdata(Broadcaster_io_ddr_in_0_bits_tdata),
    .io_ddr_in_0_bits_tkeep(Broadcaster_io_ddr_in_0_bits_tkeep),
    .io_ddr_in_0_bits_tlast(Broadcaster_io_ddr_in_0_bits_tlast),
    .io_ddr_in_1_ready(Broadcaster_io_ddr_in_1_ready),
    .io_ddr_in_1_valid(Broadcaster_io_ddr_in_1_valid),
    .io_ddr_in_1_bits_tdata(Broadcaster_io_ddr_in_1_bits_tdata),
    .io_ddr_in_1_bits_tkeep(Broadcaster_io_ddr_in_1_bits_tkeep),
    .io_ddr_in_1_bits_tlast(Broadcaster_io_ddr_in_1_bits_tlast),
    .io_ddr_in_2_ready(Broadcaster_io_ddr_in_2_ready),
    .io_ddr_in_2_valid(Broadcaster_io_ddr_in_2_valid),
    .io_ddr_in_2_bits_tdata(Broadcaster_io_ddr_in_2_bits_tdata),
    .io_ddr_in_2_bits_tkeep(Broadcaster_io_ddr_in_2_bits_tkeep),
    .io_ddr_in_2_bits_tlast(Broadcaster_io_ddr_in_2_bits_tlast),
    .io_ddr_in_3_ready(Broadcaster_io_ddr_in_3_ready),
    .io_ddr_in_3_valid(Broadcaster_io_ddr_in_3_valid),
    .io_ddr_in_3_bits_tdata(Broadcaster_io_ddr_in_3_bits_tdata),
    .io_ddr_in_3_bits_tkeep(Broadcaster_io_ddr_in_3_bits_tkeep),
    .io_ddr_in_3_bits_tlast(Broadcaster_io_ddr_in_3_bits_tlast),
    .io_pe_out_0_ready(Broadcaster_io_pe_out_0_ready),
    .io_pe_out_0_valid(Broadcaster_io_pe_out_0_valid),
    .io_pe_out_0_bits_tdata(Broadcaster_io_pe_out_0_bits_tdata),
    .io_pe_out_0_bits_tkeep(Broadcaster_io_pe_out_0_bits_tkeep),
    .io_pe_out_0_bits_tlast(Broadcaster_io_pe_out_0_bits_tlast),
    .io_pe_out_1_ready(Broadcaster_io_pe_out_1_ready),
    .io_pe_out_1_valid(Broadcaster_io_pe_out_1_valid),
    .io_pe_out_1_bits_tdata(Broadcaster_io_pe_out_1_bits_tdata),
    .io_pe_out_1_bits_tkeep(Broadcaster_io_pe_out_1_bits_tkeep),
    .io_pe_out_1_bits_tlast(Broadcaster_io_pe_out_1_bits_tlast),
    .io_pe_out_2_ready(Broadcaster_io_pe_out_2_ready),
    .io_pe_out_2_valid(Broadcaster_io_pe_out_2_valid),
    .io_pe_out_2_bits_tdata(Broadcaster_io_pe_out_2_bits_tdata),
    .io_pe_out_2_bits_tkeep(Broadcaster_io_pe_out_2_bits_tkeep),
    .io_pe_out_2_bits_tlast(Broadcaster_io_pe_out_2_bits_tlast),
    .io_pe_out_3_ready(Broadcaster_io_pe_out_3_ready),
    .io_pe_out_3_valid(Broadcaster_io_pe_out_3_valid),
    .io_pe_out_3_bits_tdata(Broadcaster_io_pe_out_3_bits_tdata),
    .io_pe_out_3_bits_tkeep(Broadcaster_io_pe_out_3_bits_tkeep),
    .io_pe_out_3_bits_tlast(Broadcaster_io_pe_out_3_bits_tlast),
    .io_pe_out_4_ready(Broadcaster_io_pe_out_4_ready),
    .io_pe_out_4_valid(Broadcaster_io_pe_out_4_valid),
    .io_pe_out_4_bits_tdata(Broadcaster_io_pe_out_4_bits_tdata),
    .io_pe_out_4_bits_tkeep(Broadcaster_io_pe_out_4_bits_tkeep),
    .io_pe_out_4_bits_tlast(Broadcaster_io_pe_out_4_bits_tlast),
    .io_pe_out_5_ready(Broadcaster_io_pe_out_5_ready),
    .io_pe_out_5_valid(Broadcaster_io_pe_out_5_valid),
    .io_pe_out_5_bits_tdata(Broadcaster_io_pe_out_5_bits_tdata),
    .io_pe_out_5_bits_tkeep(Broadcaster_io_pe_out_5_bits_tkeep),
    .io_pe_out_5_bits_tlast(Broadcaster_io_pe_out_5_bits_tlast),
    .io_pe_out_6_ready(Broadcaster_io_pe_out_6_ready),
    .io_pe_out_6_valid(Broadcaster_io_pe_out_6_valid),
    .io_pe_out_6_bits_tdata(Broadcaster_io_pe_out_6_bits_tdata),
    .io_pe_out_6_bits_tkeep(Broadcaster_io_pe_out_6_bits_tkeep),
    .io_pe_out_6_bits_tlast(Broadcaster_io_pe_out_6_bits_tlast),
    .io_pe_out_7_ready(Broadcaster_io_pe_out_7_ready),
    .io_pe_out_7_valid(Broadcaster_io_pe_out_7_valid),
    .io_pe_out_7_bits_tdata(Broadcaster_io_pe_out_7_bits_tdata),
    .io_pe_out_7_bits_tkeep(Broadcaster_io_pe_out_7_bits_tkeep),
    .io_pe_out_7_bits_tlast(Broadcaster_io_pe_out_7_bits_tlast),
    .io_pe_out_8_ready(Broadcaster_io_pe_out_8_ready),
    .io_pe_out_8_valid(Broadcaster_io_pe_out_8_valid),
    .io_pe_out_8_bits_tdata(Broadcaster_io_pe_out_8_bits_tdata),
    .io_pe_out_8_bits_tkeep(Broadcaster_io_pe_out_8_bits_tkeep),
    .io_pe_out_8_bits_tlast(Broadcaster_io_pe_out_8_bits_tlast),
    .io_pe_out_9_ready(Broadcaster_io_pe_out_9_ready),
    .io_pe_out_9_valid(Broadcaster_io_pe_out_9_valid),
    .io_pe_out_9_bits_tdata(Broadcaster_io_pe_out_9_bits_tdata),
    .io_pe_out_9_bits_tkeep(Broadcaster_io_pe_out_9_bits_tkeep),
    .io_pe_out_9_bits_tlast(Broadcaster_io_pe_out_9_bits_tlast),
    .io_pe_out_10_ready(Broadcaster_io_pe_out_10_ready),
    .io_pe_out_10_valid(Broadcaster_io_pe_out_10_valid),
    .io_pe_out_10_bits_tdata(Broadcaster_io_pe_out_10_bits_tdata),
    .io_pe_out_10_bits_tkeep(Broadcaster_io_pe_out_10_bits_tkeep),
    .io_pe_out_10_bits_tlast(Broadcaster_io_pe_out_10_bits_tlast),
    .io_pe_out_11_ready(Broadcaster_io_pe_out_11_ready),
    .io_pe_out_11_valid(Broadcaster_io_pe_out_11_valid),
    .io_pe_out_11_bits_tdata(Broadcaster_io_pe_out_11_bits_tdata),
    .io_pe_out_11_bits_tkeep(Broadcaster_io_pe_out_11_bits_tkeep),
    .io_pe_out_11_bits_tlast(Broadcaster_io_pe_out_11_bits_tlast),
    .io_pe_out_12_ready(Broadcaster_io_pe_out_12_ready),
    .io_pe_out_12_valid(Broadcaster_io_pe_out_12_valid),
    .io_pe_out_12_bits_tdata(Broadcaster_io_pe_out_12_bits_tdata),
    .io_pe_out_12_bits_tkeep(Broadcaster_io_pe_out_12_bits_tkeep),
    .io_pe_out_12_bits_tlast(Broadcaster_io_pe_out_12_bits_tlast),
    .io_pe_out_13_ready(Broadcaster_io_pe_out_13_ready),
    .io_pe_out_13_valid(Broadcaster_io_pe_out_13_valid),
    .io_pe_out_13_bits_tdata(Broadcaster_io_pe_out_13_bits_tdata),
    .io_pe_out_13_bits_tkeep(Broadcaster_io_pe_out_13_bits_tkeep),
    .io_pe_out_13_bits_tlast(Broadcaster_io_pe_out_13_bits_tlast),
    .io_pe_out_14_ready(Broadcaster_io_pe_out_14_ready),
    .io_pe_out_14_valid(Broadcaster_io_pe_out_14_valid),
    .io_pe_out_14_bits_tdata(Broadcaster_io_pe_out_14_bits_tdata),
    .io_pe_out_14_bits_tkeep(Broadcaster_io_pe_out_14_bits_tkeep),
    .io_pe_out_14_bits_tlast(Broadcaster_io_pe_out_14_bits_tlast),
    .io_pe_out_15_ready(Broadcaster_io_pe_out_15_ready),
    .io_pe_out_15_valid(Broadcaster_io_pe_out_15_valid),
    .io_pe_out_15_bits_tdata(Broadcaster_io_pe_out_15_bits_tdata),
    .io_pe_out_15_bits_tkeep(Broadcaster_io_pe_out_15_bits_tkeep),
    .io_pe_out_15_bits_tlast(Broadcaster_io_pe_out_15_bits_tlast)
  );
  assign io_config_awready = controls_io_config_awready; // @[nf_arm_doce_top_main.scala 141:22]
  assign io_config_arready = controls_io_config_arready; // @[nf_arm_doce_top_main.scala 141:22]
  assign io_config_wready = controls_io_config_wready; // @[nf_arm_doce_top_main.scala 141:22]
  assign io_config_rdata = controls_io_config_rdata; // @[nf_arm_doce_top_main.scala 141:22]
  assign io_config_rresp = 2'h0; // @[nf_arm_doce_top_main.scala 141:22]
  assign io_config_rvalid = controls_io_config_rvalid; // @[nf_arm_doce_top_main.scala 141:22]
  assign io_config_bresp = 2'h0; // @[nf_arm_doce_top_main.scala 141:22]
  assign io_config_bvalid = controls_io_config_bvalid; // @[nf_arm_doce_top_main.scala 141:22]
  assign io_PLmemory_0_aw_valid = MemController_io_ddr_out_0_aw_valid; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_aw_bits_awaddr = MemController_io_ddr_out_0_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_aw_bits_awid = 7'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_aw_bits_awlen = 8'hf; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_aw_bits_awsize = 3'h6; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_ar_valid = MemController_io_ddr_out_0_ar_valid; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_ar_bits_araddr = MemController_io_ddr_out_0_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_ar_bits_arid = 7'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_ar_bits_arlen = 8'hf; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_ar_bits_arsize = 3'h6; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_w_valid = MemController_io_ddr_out_0_w_valid; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_w_bits_wdata = MemController_io_ddr_out_0_w_bits_wdata; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_w_bits_wstrb = 64'hffffffffffffffff; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_w_bits_wlast = MemController_io_ddr_out_0_w_bits_wlast; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_r_ready = 1'h1; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_0_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_aw_bits_awid = 7'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_ar_valid = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_ar_bits_araddr = 64'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_ar_bits_arid = 7'h40; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_ar_bits_arlen = 8'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_ar_bits_arsize = 3'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_ar_bits_arburst = 2'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_w_bits_wdata = 512'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_w_bits_wstrb = 64'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_w_bits_wlast = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_r_ready = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PLmemory_1_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 87:15]
  assign io_PSmemory_0_aw_valid = LevelCache_io_axi_0_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_0_aw_bits_awaddr = LevelCache_io_axi_0_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_0_aw_bits_awid = LevelCache_io_axi_0_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_0_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_0_aw_bits_awsize = 3'h2; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_0_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_0_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_0_ar_valid = Scatters_0_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_0_ar_bits_araddr = Scatters_0_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_0_ar_bits_arid = Scatters_0_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_0_ar_bits_arlen = Scatters_0_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_0_ar_bits_arsize = Scatters_0_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_0_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_0_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_0_w_valid = LevelCache_io_axi_0_ddr_w_valid; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_0_w_bits_wdata = LevelCache_io_axi_0_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_0_w_bits_wstrb = LevelCache_io_axi_0_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_0_w_bits_wlast = 1'h1; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_0_r_ready = Scatters_0_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 100:18]
  assign io_PSmemory_0_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 93:15]
  assign io_PSmemory_1_aw_valid = LevelCache_io_axi_1_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_1_aw_bits_awaddr = LevelCache_io_axi_1_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_1_aw_bits_awid = LevelCache_io_axi_1_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_1_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_1_aw_bits_awsize = 3'h2; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_1_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_1_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_1_ar_valid = Scatters_1_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_1_ar_bits_araddr = Scatters_1_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_1_ar_bits_arid = Scatters_1_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_1_ar_bits_arlen = Scatters_1_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_1_ar_bits_arsize = Scatters_1_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_1_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_1_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_1_w_valid = LevelCache_io_axi_1_ddr_w_valid; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_1_w_bits_wdata = LevelCache_io_axi_1_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_1_w_bits_wstrb = LevelCache_io_axi_1_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_1_w_bits_wlast = 1'h1; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_1_r_ready = Scatters_1_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 100:18]
  assign io_PSmemory_1_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 93:15]
  assign io_PSmemory_2_aw_valid = LevelCache_io_axi_2_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_2_aw_bits_awaddr = LevelCache_io_axi_2_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_2_aw_bits_awid = LevelCache_io_axi_2_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_2_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_2_aw_bits_awsize = 3'h2; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_2_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_2_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_2_ar_valid = Scatters_2_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_2_ar_bits_araddr = Scatters_2_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_2_ar_bits_arid = Scatters_2_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_2_ar_bits_arlen = Scatters_2_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_2_ar_bits_arsize = Scatters_2_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_2_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_2_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_2_w_valid = LevelCache_io_axi_2_ddr_w_valid; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_2_w_bits_wdata = LevelCache_io_axi_2_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_2_w_bits_wstrb = LevelCache_io_axi_2_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_2_w_bits_wlast = 1'h1; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_2_r_ready = Scatters_2_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 100:18]
  assign io_PSmemory_2_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 93:15]
  assign io_PSmemory_3_aw_valid = LevelCache_io_axi_3_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_3_aw_bits_awaddr = LevelCache_io_axi_3_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_3_aw_bits_awid = LevelCache_io_axi_3_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_3_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_3_aw_bits_awsize = 3'h2; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_3_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_3_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 92:16]
  assign io_PSmemory_3_ar_valid = Scatters_3_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_3_ar_bits_araddr = Scatters_3_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_3_ar_bits_arid = Scatters_3_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_3_ar_bits_arlen = Scatters_3_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_3_ar_bits_arsize = Scatters_3_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_3_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_3_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 101:19]
  assign io_PSmemory_3_w_valid = LevelCache_io_axi_3_ddr_w_valid; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_3_w_bits_wdata = LevelCache_io_axi_3_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_3_w_bits_wstrb = LevelCache_io_axi_3_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_3_w_bits_wlast = 1'h1; // @[nf_arm_doce_top_main.scala 94:15]
  assign io_PSmemory_3_r_ready = Scatters_3_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 100:18]
  assign io_PSmemory_3_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 93:15]
  assign io_Re_memory_out_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 122:29]
  assign io_Re_memory_out_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_Re_memory_out_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 52:10]
  assign io_Re_memory_out_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 53:11]
  assign io_Re_memory_out_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 54:12]
  assign io_Re_memory_out_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 55:13]
  assign io_Re_memory_out_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 56:12]
  assign io_Re_memory_out_ar_valid = 1'h0; // @[nf_arm_doce_top_main.scala 124:29]
  assign io_Re_memory_out_ar_bits_araddr = 64'h0; // @[nf_arm_doce_top.scala 33:12]
  assign io_Re_memory_out_ar_bits_arid = 6'h0; // @[nf_arm_doce_top.scala 34:10]
  assign io_Re_memory_out_ar_bits_arlen = 8'h0; // @[nf_arm_doce_top.scala 35:11]
  assign io_Re_memory_out_ar_bits_arsize = 3'h0; // @[nf_arm_doce_top.scala 36:12]
  assign io_Re_memory_out_ar_bits_arburst = 2'h0; // @[nf_arm_doce_top.scala 37:13]
  assign io_Re_memory_out_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top.scala 38:12]
  assign io_Re_memory_out_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 126:28]
  assign io_Re_memory_out_w_bits_wdata = 512'h0; // @[nf_arm_doce_top.scala 66:11]
  assign io_Re_memory_out_w_bits_wstrb = 64'h0; // @[nf_arm_doce_top.scala 67:11]
  assign io_Re_memory_out_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 68:11]
  assign io_Re_memory_out_r_ready = 1'h1; // @[nf_arm_doce_top_main.scala 127:28]
  assign io_Re_memory_out_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 128:28]
  assign io_Re_memory_in_aw_ready = 1'h1; // @[nf_arm_doce_top_main.scala 119:28]
  assign io_Re_memory_in_ar_ready = 1'h1; // @[nf_arm_doce_top_main.scala 118:28]
  assign io_Re_memory_in_w_ready = 1'h1; // @[nf_arm_doce_top_main.scala 120:27]
  assign io_Re_memory_in_r_valid = 1'h0; // @[nf_arm_doce_top_main.scala 115:27]
  assign io_Re_memory_in_r_bits_rdata = 512'h0; // @[nf_arm_doce_top.scala 88:11]
  assign io_Re_memory_in_r_bits_rid = 10'h0; // @[nf_arm_doce_top.scala 89:9]
  assign io_Re_memory_in_r_bits_rlast = 1'h0; // @[nf_arm_doce_top.scala 90:11]
  assign io_Re_memory_in_b_valid = 1'h0; // @[nf_arm_doce_top_main.scala 117:27]
  assign io_Re_memory_in_b_bits_bresp = 2'h0; // @[nf_arm_doce_top.scala 77:11]
  assign io_Re_memory_in_b_bits_bid = 10'h0; // @[nf_arm_doce_top.scala 78:9]
  assign controls_clock = clock;
  assign controls_reset = reset;
  assign controls_io_fin_0 = Applys_0_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_1 = Applys_1_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_2 = Applys_2_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_3 = Applys_3_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_4 = Applys_4_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_5 = Applys_5_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_6 = Applys_6_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_7 = Applys_7_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_8 = Applys_8_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_9 = Applys_9_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_10 = Applys_10_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_11 = Applys_11_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_12 = Applys_12_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_13 = Applys_13_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_14 = Applys_14_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_fin_15 = Applys_15_io_end; // @[nf_arm_doce_top_main.scala 109:26]
  assign controls_io_unvisited_size = MemController_io_unvisited_size; // @[nf_arm_doce_top_main.scala 143:30]
  assign controls_io_traveled_edges = _controls_io_traveled_edges_T_3 + Scatters_3_io_traveled_edges; // @[nf_arm_doce_top_main.scala 142:80]
  assign controls_io_config_awaddr = io_config_awaddr; // @[nf_arm_doce_top_main.scala 141:22]
  assign controls_io_config_awvalid = io_config_awvalid; // @[nf_arm_doce_top_main.scala 141:22]
  assign controls_io_config_araddr = io_config_araddr; // @[nf_arm_doce_top_main.scala 141:22]
  assign controls_io_config_arvalid = io_config_arvalid; // @[nf_arm_doce_top_main.scala 141:22]
  assign controls_io_config_wdata = io_config_wdata; // @[nf_arm_doce_top_main.scala 141:22]
  assign controls_io_config_wvalid = io_config_wvalid; // @[nf_arm_doce_top_main.scala 141:22]
  assign controls_io_config_rready = io_config_rready; // @[nf_arm_doce_top_main.scala 141:22]
  assign controls_io_config_bready = io_config_bready; // @[nf_arm_doce_top_main.scala 141:22]
  assign controls_io_flush_cache_end = LevelCache_io_end; // @[nf_arm_doce_top_main.scala 144:31]
  assign controls_io_signal_ack = MemController_io_signal_ack; // @[nf_arm_doce_top_main.scala 145:26]
  assign MemController_clock = clock;
  assign MemController_reset = reset;
  assign MemController_io_cacheable_out_ready = Gathers_io_ddr_in_ready; // @[nf_arm_doce_top_main.scala 88:21]
  assign MemController_io_cacheable_in_0_valid = Applys_0_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_0_bits_tdata = Applys_0_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_1_valid = Applys_1_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_1_bits_tdata = Applys_1_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_2_valid = Applys_2_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_2_bits_tdata = Applys_2_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_3_valid = Applys_3_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_3_bits_tdata = Applys_3_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_4_valid = Applys_4_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_4_bits_tdata = Applys_4_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_5_valid = Applys_5_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_5_bits_tdata = Applys_5_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_6_valid = Applys_6_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_6_bits_tdata = Applys_6_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_7_valid = Applys_7_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_7_bits_tdata = Applys_7_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_8_valid = Applys_8_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_8_bits_tdata = Applys_8_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_9_valid = Applys_9_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_9_bits_tdata = Applys_9_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_10_valid = Applys_10_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_10_bits_tdata = Applys_10_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_11_valid = Applys_11_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_11_bits_tdata = Applys_11_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_12_valid = Applys_12_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_12_bits_tdata = Applys_12_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_13_valid = Applys_13_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_13_bits_tdata = Applys_13_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_14_valid = Applys_14_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_14_bits_tdata = Applys_14_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_15_valid = Applys_15_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_cacheable_in_15_bits_tdata = Applys_15_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 108:21]
  assign MemController_io_ddr_out_0_aw_ready = io_PLmemory_0_aw_ready; // @[nf_arm_doce_top_main.scala 87:15]
  assign MemController_io_ddr_out_0_ar_ready = io_PLmemory_0_ar_ready; // @[nf_arm_doce_top_main.scala 87:15]
  assign MemController_io_ddr_out_0_w_ready = io_PLmemory_0_w_ready; // @[nf_arm_doce_top_main.scala 87:15]
  assign MemController_io_ddr_out_0_r_valid = io_PLmemory_0_r_valid; // @[nf_arm_doce_top_main.scala 87:15]
  assign MemController_io_ddr_out_0_r_bits_rdata = io_PLmemory_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 87:15]
  assign MemController_io_ddr_out_0_r_bits_rlast = io_PLmemory_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 87:15]
  assign MemController_io_tiers_base_addr_0 = {controls_io_data_9,controls_io_data_8}; // @[Cat.scala 30:58]
  assign MemController_io_tiers_base_addr_1 = {controls_io_data_11,controls_io_data_10}; // @[Cat.scala 30:58]
  assign MemController_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 168:26]
  assign MemController_io_signal = controls_io_signal & controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 167:49]
  assign MemController_io_end = controls_io_data_0[1]; // @[nf_arm_doce_top_main.scala 169:46]
  assign Applys_0_clock = clock;
  assign Applys_0_reset = reset;
  assign Applys_0_io_xbar_in_valid = Broadcaster_io_pe_out_0_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_0_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_0_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_0_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_0_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_0_io_ddr_out_ready = MemController_io_cacheable_in_0_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_1_clock = clock;
  assign Applys_1_reset = reset;
  assign Applys_1_io_xbar_in_valid = Broadcaster_io_pe_out_1_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_1_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_1_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_1_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_1_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_1_io_ddr_out_ready = MemController_io_cacheable_in_1_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_2_clock = clock;
  assign Applys_2_reset = reset;
  assign Applys_2_io_xbar_in_valid = Broadcaster_io_pe_out_2_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_2_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_2_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_2_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_2_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_2_io_ddr_out_ready = MemController_io_cacheable_in_2_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_3_clock = clock;
  assign Applys_3_reset = reset;
  assign Applys_3_io_xbar_in_valid = Broadcaster_io_pe_out_3_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_3_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_3_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_3_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_3_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_3_io_ddr_out_ready = MemController_io_cacheable_in_3_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_4_clock = clock;
  assign Applys_4_reset = reset;
  assign Applys_4_io_xbar_in_valid = Broadcaster_io_pe_out_4_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_4_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_4_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_4_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_4_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_4_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_4_io_ddr_out_ready = MemController_io_cacheable_in_4_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_5_clock = clock;
  assign Applys_5_reset = reset;
  assign Applys_5_io_xbar_in_valid = Broadcaster_io_pe_out_5_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_5_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_5_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_5_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_5_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_5_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_5_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_5_io_ddr_out_ready = MemController_io_cacheable_in_5_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_6_clock = clock;
  assign Applys_6_reset = reset;
  assign Applys_6_io_xbar_in_valid = Broadcaster_io_pe_out_6_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_6_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_6_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_6_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_6_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_6_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_6_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_6_io_ddr_out_ready = MemController_io_cacheable_in_6_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_7_clock = clock;
  assign Applys_7_reset = reset;
  assign Applys_7_io_xbar_in_valid = Broadcaster_io_pe_out_7_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_7_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_7_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_7_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_7_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_7_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_7_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_7_io_ddr_out_ready = MemController_io_cacheable_in_7_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_8_clock = clock;
  assign Applys_8_reset = reset;
  assign Applys_8_io_xbar_in_valid = Broadcaster_io_pe_out_8_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_8_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_8_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_8_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_8_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_8_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_8_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_8_io_ddr_out_ready = MemController_io_cacheable_in_8_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_9_clock = clock;
  assign Applys_9_reset = reset;
  assign Applys_9_io_xbar_in_valid = Broadcaster_io_pe_out_9_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_9_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_9_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_9_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_9_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_9_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_9_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_9_io_ddr_out_ready = MemController_io_cacheable_in_9_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_10_clock = clock;
  assign Applys_10_reset = reset;
  assign Applys_10_io_xbar_in_valid = Broadcaster_io_pe_out_10_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_10_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_10_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_10_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_10_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_10_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_10_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_10_io_ddr_out_ready = MemController_io_cacheable_in_10_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_11_clock = clock;
  assign Applys_11_reset = reset;
  assign Applys_11_io_xbar_in_valid = Broadcaster_io_pe_out_11_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_11_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_11_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_11_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_11_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_11_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_11_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_11_io_ddr_out_ready = MemController_io_cacheable_in_11_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_12_clock = clock;
  assign Applys_12_reset = reset;
  assign Applys_12_io_xbar_in_valid = Broadcaster_io_pe_out_12_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_12_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_12_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_12_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_12_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_12_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_12_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_12_io_ddr_out_ready = MemController_io_cacheable_in_12_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_13_clock = clock;
  assign Applys_13_reset = reset;
  assign Applys_13_io_xbar_in_valid = Broadcaster_io_pe_out_13_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_13_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_13_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_13_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_13_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_13_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_13_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_13_io_ddr_out_ready = MemController_io_cacheable_in_13_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_14_clock = clock;
  assign Applys_14_reset = reset;
  assign Applys_14_io_xbar_in_valid = Broadcaster_io_pe_out_14_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_14_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_14_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_14_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_14_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_14_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_14_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_14_io_ddr_out_ready = MemController_io_cacheable_in_14_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Applys_15_clock = clock;
  assign Applys_15_reset = reset;
  assign Applys_15_io_xbar_in_valid = Broadcaster_io_pe_out_15_valid; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_15_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_15_bits_tdata; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_15_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_15_bits_tkeep; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_15_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_15_bits_tlast; // @[nf_arm_doce_top_main.scala 107:21]
  assign Applys_15_io_ddr_out_ready = MemController_io_cacheable_in_15_ready; // @[nf_arm_doce_top_main.scala 108:21]
  assign Gathers_clock = clock;
  assign Gathers_reset = reset;
  assign Gathers_io_ddr_in_valid = MemController_io_cacheable_out_valid; // @[nf_arm_doce_top_main.scala 88:21]
  assign Gathers_io_ddr_in_bits_tdata = MemController_io_cacheable_out_bits_tdata; // @[nf_arm_doce_top_main.scala 88:21]
  assign Gathers_io_ddr_in_bits_tkeep = MemController_io_cacheable_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 88:21]
  assign Gathers_io_gather_out_0_ready = Scatters_0_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 99:22]
  assign Gathers_io_gather_out_1_ready = Scatters_1_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 99:22]
  assign Gathers_io_gather_out_2_ready = Scatters_2_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 99:22]
  assign Gathers_io_gather_out_3_ready = Scatters_3_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 99:22]
  assign Gathers_io_level_cache_out_ready = LevelCache_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 89:27]
  assign LevelCache_clock = clock;
  assign LevelCache_reset = reset;
  assign LevelCache_io_axi_0_ddr_aw_ready = io_PSmemory_0_aw_ready; // @[nf_arm_doce_top_main.scala 92:16]
  assign LevelCache_io_axi_0_ddr_w_ready = io_PSmemory_0_w_ready; // @[nf_arm_doce_top_main.scala 94:15]
  assign LevelCache_io_axi_1_ddr_aw_ready = io_PSmemory_1_aw_ready; // @[nf_arm_doce_top_main.scala 92:16]
  assign LevelCache_io_axi_1_ddr_w_ready = io_PSmemory_1_w_ready; // @[nf_arm_doce_top_main.scala 94:15]
  assign LevelCache_io_axi_2_ddr_aw_ready = io_PSmemory_2_aw_ready; // @[nf_arm_doce_top_main.scala 92:16]
  assign LevelCache_io_axi_2_ddr_w_ready = io_PSmemory_2_w_ready; // @[nf_arm_doce_top_main.scala 94:15]
  assign LevelCache_io_axi_3_ddr_aw_ready = io_PSmemory_3_aw_ready; // @[nf_arm_doce_top_main.scala 92:16]
  assign LevelCache_io_axi_3_ddr_w_ready = io_PSmemory_3_w_ready; // @[nf_arm_doce_top_main.scala 94:15]
  assign LevelCache_io_gather_in_valid = Gathers_io_level_cache_out_valid; // @[nf_arm_doce_top_main.scala 89:27]
  assign LevelCache_io_gather_in_bits_tdata = Gathers_io_level_cache_out_bits_tdata; // @[nf_arm_doce_top_main.scala 89:27]
  assign LevelCache_io_gather_in_bits_tkeep = {{48'd0}, Gathers_io_level_cache_out_bits_tkeep}; // @[nf_arm_doce_top_main.scala 89:27]
  assign LevelCache_io_gather_in_bits_tlast = Gathers_io_level_cache_out_bits_tlast; // @[nf_arm_doce_top_main.scala 89:27]
  assign LevelCache_io_level = controls_io_level; // @[nf_arm_doce_top_main.scala 150:23]
  assign LevelCache_io_level_base_addr = {controls_io_data_6,controls_io_data_5}; // @[Cat.scala 30:58]
  assign LevelCache_io_flush = controls_io_flush_cache; // @[nf_arm_doce_top_main.scala 148:23]
  assign Scatters_0_clock = clock;
  assign Scatters_0_reset = reset;
  assign Scatters_0_io_ddr_ar_ready = io_PSmemory_0_ar_ready; // @[nf_arm_doce_top_main.scala 101:19]
  assign Scatters_0_io_ddr_r_valid = io_PSmemory_0_r_valid; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_0_io_ddr_r_bits_rdata = io_PSmemory_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_0_io_ddr_r_bits_rid = io_PSmemory_0_r_bits_rid; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_0_io_ddr_r_bits_rlast = io_PSmemory_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_0_io_gather_in_valid = Gathers_io_gather_out_0_valid; // @[nf_arm_doce_top_main.scala 99:22]
  assign Scatters_0_io_gather_in_bits_tdata = Gathers_io_gather_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 99:22]
  assign Scatters_0_io_xbar_out_ready = Broadcaster_io_ddr_in_0_ready; // @[nf_arm_doce_top_main.scala 102:32]
  assign Scatters_0_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_0_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_0_io_signal = controls_io_signal & controls_io_signal_ack | controls_io_start; // @[nf_arm_doce_top_main.scala 154:69]
  assign Scatters_0_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 158:20]
  assign Scatters_0_io_root = controls_io_data_7; // @[nf_arm_doce_top_main.scala 153:17]
  assign Scatters_0_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 162:75]
  assign Scatters_1_clock = clock;
  assign Scatters_1_reset = reset;
  assign Scatters_1_io_ddr_ar_ready = io_PSmemory_1_ar_ready; // @[nf_arm_doce_top_main.scala 101:19]
  assign Scatters_1_io_ddr_r_valid = io_PSmemory_1_r_valid; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_1_io_ddr_r_bits_rdata = io_PSmemory_1_r_bits_rdata; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_1_io_ddr_r_bits_rid = io_PSmemory_1_r_bits_rid; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_1_io_ddr_r_bits_rlast = io_PSmemory_1_r_bits_rlast; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_1_io_gather_in_valid = Gathers_io_gather_out_1_valid; // @[nf_arm_doce_top_main.scala 99:22]
  assign Scatters_1_io_gather_in_bits_tdata = Gathers_io_gather_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 99:22]
  assign Scatters_1_io_xbar_out_ready = Broadcaster_io_ddr_in_1_ready; // @[nf_arm_doce_top_main.scala 102:32]
  assign Scatters_1_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_1_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_1_io_signal = controls_io_signal & controls_io_signal_ack | controls_io_start; // @[nf_arm_doce_top_main.scala 154:69]
  assign Scatters_1_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 162:75]
  assign Scatters_2_clock = clock;
  assign Scatters_2_reset = reset;
  assign Scatters_2_io_ddr_ar_ready = io_PSmemory_2_ar_ready; // @[nf_arm_doce_top_main.scala 101:19]
  assign Scatters_2_io_ddr_r_valid = io_PSmemory_2_r_valid; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_2_io_ddr_r_bits_rdata = io_PSmemory_2_r_bits_rdata; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_2_io_ddr_r_bits_rid = io_PSmemory_2_r_bits_rid; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_2_io_ddr_r_bits_rlast = io_PSmemory_2_r_bits_rlast; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_2_io_gather_in_valid = Gathers_io_gather_out_2_valid; // @[nf_arm_doce_top_main.scala 99:22]
  assign Scatters_2_io_gather_in_bits_tdata = Gathers_io_gather_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 99:22]
  assign Scatters_2_io_xbar_out_ready = Broadcaster_io_ddr_in_2_ready; // @[nf_arm_doce_top_main.scala 102:32]
  assign Scatters_2_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_2_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_2_io_signal = controls_io_signal & controls_io_signal_ack | controls_io_start; // @[nf_arm_doce_top_main.scala 154:69]
  assign Scatters_2_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 162:75]
  assign Scatters_3_clock = clock;
  assign Scatters_3_reset = reset;
  assign Scatters_3_io_ddr_ar_ready = io_PSmemory_3_ar_ready; // @[nf_arm_doce_top_main.scala 101:19]
  assign Scatters_3_io_ddr_r_valid = io_PSmemory_3_r_valid; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_3_io_ddr_r_bits_rdata = io_PSmemory_3_r_bits_rdata; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_3_io_ddr_r_bits_rid = io_PSmemory_3_r_bits_rid; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_3_io_ddr_r_bits_rlast = io_PSmemory_3_r_bits_rlast; // @[nf_arm_doce_top_main.scala 100:18]
  assign Scatters_3_io_gather_in_valid = Gathers_io_gather_out_3_valid; // @[nf_arm_doce_top_main.scala 99:22]
  assign Scatters_3_io_gather_in_bits_tdata = Gathers_io_gather_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 99:22]
  assign Scatters_3_io_xbar_out_ready = Broadcaster_io_ddr_in_3_ready; // @[nf_arm_doce_top_main.scala 102:32]
  assign Scatters_3_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_3_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_3_io_signal = controls_io_signal & controls_io_signal_ack | controls_io_start; // @[nf_arm_doce_top_main.scala 154:69]
  assign Scatters_3_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 162:75]
  assign Broadcaster_clock = clock;
  assign Broadcaster_reset = reset;
  assign Broadcaster_io_ddr_in_0_valid = Scatters_0_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_0_bits_tdata = Scatters_0_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_0_bits_tkeep = Scatters_0_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_0_bits_tlast = Scatters_0_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_1_valid = Scatters_1_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_1_bits_tdata = Scatters_1_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_1_bits_tkeep = Scatters_1_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_1_bits_tlast = Scatters_1_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_2_valid = Scatters_2_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_2_bits_tdata = Scatters_2_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_2_bits_tkeep = Scatters_2_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_2_bits_tlast = Scatters_2_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_3_valid = Scatters_3_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_3_bits_tdata = Scatters_3_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_3_bits_tkeep = Scatters_3_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_ddr_in_3_bits_tlast = Scatters_3_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 102:32]
  assign Broadcaster_io_pe_out_0_ready = Applys_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_1_ready = Applys_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_2_ready = Applys_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_3_ready = Applys_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_4_ready = Applys_4_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_5_ready = Applys_5_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_6_ready = Applys_6_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_7_ready = Applys_7_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_8_ready = Applys_8_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_9_ready = Applys_9_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_10_ready = Applys_10_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_11_ready = Applys_11_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_12_ready = Applys_12_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_13_ready = Applys_13_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_14_ready = Applys_14_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  assign Broadcaster_io_pe_out_15_ready = Applys_15_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 107:21]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      ar_ready_counter1 <= 31'h0; // @[Counter.scala 60:40]
    end else if (_T_5) begin // @[Counter.scala 118:17]
      if (wrap_wrap) begin // @[Counter.scala 86:20]
        ar_ready_counter1 <= 31'h0; // @[Counter.scala 86:28]
      end else begin
        ar_ready_counter1 <= _wrap_value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[nf_arm_doce_top_main.scala 49:34]
      axi_ready_counter_0 <= 32'h0; // @[nf_arm_doce_top_main.scala 49:34]
    end else if (_T_14) begin // @[nf_arm_doce_top_main.scala 55:43]
      axi_ready_counter_0 <= _axi_ready_counter_0_T_1; // @[nf_arm_doce_top_main.scala 56:10]
    end
    if (reset) begin // @[nf_arm_doce_top_main.scala 49:34]
      axi_ready_counter_1 <= 32'h0; // @[nf_arm_doce_top_main.scala 49:34]
    end else if (_T_23) begin // @[nf_arm_doce_top_main.scala 55:43]
      axi_ready_counter_1 <= _axi_ready_counter_1_T_1; // @[nf_arm_doce_top_main.scala 56:10]
    end
    if (reset) begin // @[nf_arm_doce_top_main.scala 49:34]
      axi_ready_counter_2 <= 32'h0; // @[nf_arm_doce_top_main.scala 49:34]
    end else if (_T_32) begin // @[nf_arm_doce_top_main.scala 55:43]
      axi_ready_counter_2 <= _axi_ready_counter_2_T_1; // @[nf_arm_doce_top_main.scala 56:10]
    end
    if (reset) begin // @[nf_arm_doce_top_main.scala 49:34]
      axi_ready_counter_3 <= 32'h0; // @[nf_arm_doce_top_main.scala 49:34]
    end else if (_T_41) begin // @[nf_arm_doce_top_main.scala 55:43]
      axi_ready_counter_3 <= _axi_ready_counter_3_T_1; // @[nf_arm_doce_top_main.scala 56:10]
    end
    if (reset) begin // @[nf_arm_doce_top_main.scala 60:38]
      axi_all_ready_counter <= 32'h0; // @[nf_arm_doce_top_main.scala 60:38]
    end else if (_T_74) begin // @[nf_arm_doce_top_main.scala 70:40]
      axi_all_ready_counter <= _axi_all_ready_counter_T_1; // @[nf_arm_doce_top_main.scala 71:27]
    end
    if (reset) begin // @[nf_arm_doce_top_main.scala 73:40]
      axi_r_all_ready_counter <= 32'h0; // @[nf_arm_doce_top_main.scala 73:40]
    end else if (_T_91) begin // @[nf_arm_doce_top_main.scala 83:40]
      axi_r_all_ready_counter <= _axi_r_all_ready_counter_T_1; // @[nf_arm_doce_top_main.scala 84:29]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ar_ready_counter1 = _RAND_0[30:0];
  _RAND_1 = {1{`RANDOM}};
  axi_ready_counter_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  axi_ready_counter_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  axi_ready_counter_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  axi_ready_counter_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  axi_all_ready_counter = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  axi_r_all_ready_counter = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
