module LookupTable(
  input         clock,
  input         reset,
  output [31:0] io_data_0,
  output [31:0] io_data_1,
  output [31:0] io_data_2,
  output [31:0] io_data_3,
  output [31:0] io_data_4,
  output [31:0] io_data_7,
  output [31:0] io_data_12,
  output [31:0] io_data_13,
  output [31:0] io_data_16,
  output [31:0] io_data_17,
  output [31:0] io_data_18,
  output [31:0] io_data_19,
  output [31:0] io_data_20,
  output [31:0] io_data_21,
  output [31:0] io_data_22,
  output [31:0] io_data_23,
  output [31:0] io_data_24,
  output [31:0] io_data_25,
  output [31:0] io_data_26,
  output [31:0] io_data_27,
  output [31:0] io_data_28,
  output [31:0] io_data_29,
  input  [31:0] io_dataIn_0,
  input  [31:0] io_dataIn_1,
  input         io_writeFlag_0,
  input         io_writeFlag_1,
  input  [4:0]  io_wptr_0,
  input  [4:0]  io_wptr_1,
  input  [63:0] config_awaddr,
  input         config_awvalid,
  output        config_awready,
  input  [63:0] config_araddr,
  input         config_arvalid,
  output        config_arready,
  input  [31:0] config_wdata,
  input         config_wvalid,
  output        config_wready,
  output [31:0] config_rdata,
  output        config_rvalid,
  input         config_rready,
  output        config_bvalid,
  input         config_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] table_0; // @[util.scala 16:22]
  reg [31:0] table_1; // @[util.scala 16:22]
  reg [31:0] table_2; // @[util.scala 16:22]
  reg [31:0] table_3; // @[util.scala 16:22]
  reg [31:0] table_4; // @[util.scala 16:22]
  reg [31:0] table_5; // @[util.scala 16:22]
  reg [31:0] table_6; // @[util.scala 16:22]
  reg [31:0] table_7; // @[util.scala 16:22]
  reg [31:0] table_8; // @[util.scala 16:22]
  reg [31:0] table_9; // @[util.scala 16:22]
  reg [31:0] table_10; // @[util.scala 16:22]
  reg [31:0] table_11; // @[util.scala 16:22]
  reg [31:0] table_12; // @[util.scala 16:22]
  (*dont_touch = "true" *)reg [31:0] table_13; // @[util.scala 16:22]
  reg [31:0] table_14; // @[util.scala 16:22]
  reg [31:0] table_15; // @[util.scala 16:22]
  reg [31:0] table_16; // @[util.scala 16:22]
  reg [31:0] table_17; // @[util.scala 16:22]
  reg [31:0] table_18; // @[util.scala 16:22]
  reg [31:0] table_19; // @[util.scala 16:22]
  reg [31:0] table_20; // @[util.scala 16:22]
  reg [31:0] table_21; // @[util.scala 16:22]
  reg [31:0] table_22; // @[util.scala 16:22]
  reg [31:0] table_23; // @[util.scala 16:22]
  reg [31:0] table_24; // @[util.scala 16:22]
  reg [31:0] table_25; // @[util.scala 16:22]
  reg [31:0] table_26; // @[util.scala 16:22]
  reg [31:0] table_27; // @[util.scala 16:22]
  reg [31:0] table_28; // @[util.scala 16:22]
  reg [31:0] table_29; // @[util.scala 16:22]
  reg [31:0] table_30; // @[util.scala 16:22]
  reg [31:0] table_31; // @[util.scala 16:22]
  reg [2:0] status; // @[util.scala 26:23]
  wire [2:0] _GEN_3 = config_bready ? 3'h0 : status; // @[util.scala 41:24 util.scala 42:14 util.scala 26:23]
  wire [2:0] _GEN_4 = config_rready ? 3'h0 : status; // @[util.scala 47:25 util.scala 48:14 util.scala 26:23]
  wire [2:0] _GEN_5 = status == 3'h5 ? _GEN_4 : status; // @[util.scala 46:36 util.scala 26:23]
  wire [2:0] _GEN_6 = status == 3'h4 ? 3'h5 : _GEN_5; // @[util.scala 44:35 util.scala 45:12]
  wire [2:0] _GEN_7 = status == 3'h3 ? _GEN_3 : _GEN_6; // @[util.scala 40:35]
  wire  wvalid = config_wvalid & config_wready; // @[util.scala 64:30]
  reg [4:0] ewaddr; // @[util.scala 65:19]
  wire  _T_7 = io_writeFlag_0 & io_writeFlag_1; // @[util.scala 70:39]
  wire [31:0] _GEN_12 = 5'h0 == ewaddr ? config_wdata : table_0; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_13 = 5'h1 == ewaddr ? config_wdata : table_1; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_14 = 5'h2 == ewaddr ? config_wdata : table_2; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_15 = 5'h3 == ewaddr ? config_wdata : table_3; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_16 = 5'h4 == ewaddr ? config_wdata : table_4; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_17 = 5'h5 == ewaddr ? config_wdata : table_5; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_18 = 5'h6 == ewaddr ? config_wdata : table_6; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_19 = 5'h7 == ewaddr ? config_wdata : table_7; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_20 = 5'h8 == ewaddr ? config_wdata : table_8; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_21 = 5'h9 == ewaddr ? config_wdata : table_9; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_22 = 5'ha == ewaddr ? config_wdata : table_10; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_23 = 5'hb == ewaddr ? config_wdata : table_11; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_24 = 5'hc == ewaddr ? config_wdata : table_12; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_25 = 5'hd == ewaddr ? config_wdata : table_13; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_26 = 5'he == ewaddr ? config_wdata : table_14; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_27 = 5'hf == ewaddr ? config_wdata : table_15; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_28 = 5'h10 == ewaddr ? config_wdata : table_16; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_29 = 5'h11 == ewaddr ? config_wdata : table_17; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_30 = 5'h12 == ewaddr ? config_wdata : table_18; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_31 = 5'h13 == ewaddr ? config_wdata : table_19; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_32 = 5'h14 == ewaddr ? config_wdata : table_20; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_33 = 5'h15 == ewaddr ? config_wdata : table_21; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_34 = 5'h16 == ewaddr ? config_wdata : table_22; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_35 = 5'h17 == ewaddr ? config_wdata : table_23; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_36 = 5'h18 == ewaddr ? config_wdata : table_24; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_37 = 5'h19 == ewaddr ? config_wdata : table_25; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_38 = 5'h1a == ewaddr ? config_wdata : table_26; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_39 = 5'h1b == ewaddr ? config_wdata : table_27; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_40 = 5'h1c == ewaddr ? config_wdata : table_28; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_41 = 5'h1d == ewaddr ? config_wdata : table_29; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_42 = 5'h1e == ewaddr ? config_wdata : table_30; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_43 = 5'h1f == ewaddr ? config_wdata : table_31; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_44 = 5'h0 == io_wptr_0 ? io_dataIn_0 : _GEN_12; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_45 = 5'h1 == io_wptr_0 ? io_dataIn_0 : _GEN_13; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_46 = 5'h2 == io_wptr_0 ? io_dataIn_0 : _GEN_14; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_47 = 5'h3 == io_wptr_0 ? io_dataIn_0 : _GEN_15; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_48 = 5'h4 == io_wptr_0 ? io_dataIn_0 : _GEN_16; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_49 = 5'h5 == io_wptr_0 ? io_dataIn_0 : _GEN_17; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_50 = 5'h6 == io_wptr_0 ? io_dataIn_0 : _GEN_18; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_51 = 5'h7 == io_wptr_0 ? io_dataIn_0 : _GEN_19; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_52 = 5'h8 == io_wptr_0 ? io_dataIn_0 : _GEN_20; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_53 = 5'h9 == io_wptr_0 ? io_dataIn_0 : _GEN_21; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_54 = 5'ha == io_wptr_0 ? io_dataIn_0 : _GEN_22; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_55 = 5'hb == io_wptr_0 ? io_dataIn_0 : _GEN_23; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_56 = 5'hc == io_wptr_0 ? io_dataIn_0 : _GEN_24; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_57 = 5'hd == io_wptr_0 ? io_dataIn_0 : _GEN_25; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_58 = 5'he == io_wptr_0 ? io_dataIn_0 : _GEN_26; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_59 = 5'hf == io_wptr_0 ? io_dataIn_0 : _GEN_27; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_60 = 5'h10 == io_wptr_0 ? io_dataIn_0 : _GEN_28; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_61 = 5'h11 == io_wptr_0 ? io_dataIn_0 : _GEN_29; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_62 = 5'h12 == io_wptr_0 ? io_dataIn_0 : _GEN_30; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_63 = 5'h13 == io_wptr_0 ? io_dataIn_0 : _GEN_31; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_64 = 5'h14 == io_wptr_0 ? io_dataIn_0 : _GEN_32; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_65 = 5'h15 == io_wptr_0 ? io_dataIn_0 : _GEN_33; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_66 = 5'h16 == io_wptr_0 ? io_dataIn_0 : _GEN_34; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_67 = 5'h17 == io_wptr_0 ? io_dataIn_0 : _GEN_35; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_68 = 5'h18 == io_wptr_0 ? io_dataIn_0 : _GEN_36; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_69 = 5'h19 == io_wptr_0 ? io_dataIn_0 : _GEN_37; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_70 = 5'h1a == io_wptr_0 ? io_dataIn_0 : _GEN_38; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_71 = 5'h1b == io_wptr_0 ? io_dataIn_0 : _GEN_39; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_72 = 5'h1c == io_wptr_0 ? io_dataIn_0 : _GEN_40; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_73 = 5'h1d == io_wptr_0 ? io_dataIn_0 : _GEN_41; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_74 = 5'h1e == io_wptr_0 ? io_dataIn_0 : _GEN_42; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_75 = 5'h1f == io_wptr_0 ? io_dataIn_0 : _GEN_43; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_204 = 5'h0 == io_wptr_1 ? io_dataIn_1 : _GEN_12; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_205 = 5'h1 == io_wptr_1 ? io_dataIn_1 : _GEN_13; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_206 = 5'h2 == io_wptr_1 ? io_dataIn_1 : _GEN_14; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_207 = 5'h3 == io_wptr_1 ? io_dataIn_1 : _GEN_15; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_208 = 5'h4 == io_wptr_1 ? io_dataIn_1 : _GEN_16; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_209 = 5'h5 == io_wptr_1 ? io_dataIn_1 : _GEN_17; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_210 = 5'h6 == io_wptr_1 ? io_dataIn_1 : _GEN_18; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_211 = 5'h7 == io_wptr_1 ? io_dataIn_1 : _GEN_19; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_212 = 5'h8 == io_wptr_1 ? io_dataIn_1 : _GEN_20; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_213 = 5'h9 == io_wptr_1 ? io_dataIn_1 : _GEN_21; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_214 = 5'ha == io_wptr_1 ? io_dataIn_1 : _GEN_22; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_215 = 5'hb == io_wptr_1 ? io_dataIn_1 : _GEN_23; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_216 = 5'hc == io_wptr_1 ? io_dataIn_1 : _GEN_24; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_217 = 5'hd == io_wptr_1 ? io_dataIn_1 : _GEN_25; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_218 = 5'he == io_wptr_1 ? io_dataIn_1 : _GEN_26; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_219 = 5'hf == io_wptr_1 ? io_dataIn_1 : _GEN_27; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_220 = 5'h10 == io_wptr_1 ? io_dataIn_1 : _GEN_28; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_221 = 5'h11 == io_wptr_1 ? io_dataIn_1 : _GEN_29; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_222 = 5'h12 == io_wptr_1 ? io_dataIn_1 : _GEN_30; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_223 = 5'h13 == io_wptr_1 ? io_dataIn_1 : _GEN_31; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_224 = 5'h14 == io_wptr_1 ? io_dataIn_1 : _GEN_32; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_225 = 5'h15 == io_wptr_1 ? io_dataIn_1 : _GEN_33; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_226 = 5'h16 == io_wptr_1 ? io_dataIn_1 : _GEN_34; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_227 = 5'h17 == io_wptr_1 ? io_dataIn_1 : _GEN_35; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_228 = 5'h18 == io_wptr_1 ? io_dataIn_1 : _GEN_36; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_229 = 5'h19 == io_wptr_1 ? io_dataIn_1 : _GEN_37; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_230 = 5'h1a == io_wptr_1 ? io_dataIn_1 : _GEN_38; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_231 = 5'h1b == io_wptr_1 ? io_dataIn_1 : _GEN_39; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_232 = 5'h1c == io_wptr_1 ? io_dataIn_1 : _GEN_40; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_233 = 5'h1d == io_wptr_1 ? io_dataIn_1 : _GEN_41; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_234 = 5'h1e == io_wptr_1 ? io_dataIn_1 : _GEN_42; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_235 = 5'h1f == io_wptr_1 ? io_dataIn_1 : _GEN_43; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_268 = 5'h0 == io_wptr_0 ? io_dataIn_0 : table_0; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_269 = 5'h1 == io_wptr_0 ? io_dataIn_0 : table_1; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_270 = 5'h2 == io_wptr_0 ? io_dataIn_0 : table_2; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_271 = 5'h3 == io_wptr_0 ? io_dataIn_0 : table_3; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_272 = 5'h4 == io_wptr_0 ? io_dataIn_0 : table_4; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_273 = 5'h5 == io_wptr_0 ? io_dataIn_0 : table_5; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_274 = 5'h6 == io_wptr_0 ? io_dataIn_0 : table_6; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_275 = 5'h7 == io_wptr_0 ? io_dataIn_0 : table_7; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_276 = 5'h8 == io_wptr_0 ? io_dataIn_0 : table_8; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_277 = 5'h9 == io_wptr_0 ? io_dataIn_0 : table_9; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_278 = 5'ha == io_wptr_0 ? io_dataIn_0 : table_10; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_279 = 5'hb == io_wptr_0 ? io_dataIn_0 : table_11; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_280 = 5'hc == io_wptr_0 ? io_dataIn_0 : table_12; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_281 = 5'hd == io_wptr_0 ? io_dataIn_0 : table_13; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_282 = 5'he == io_wptr_0 ? io_dataIn_0 : table_14; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_283 = 5'hf == io_wptr_0 ? io_dataIn_0 : table_15; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_284 = 5'h10 == io_wptr_0 ? io_dataIn_0 : table_16; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_285 = 5'h11 == io_wptr_0 ? io_dataIn_0 : table_17; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_286 = 5'h12 == io_wptr_0 ? io_dataIn_0 : table_18; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_287 = 5'h13 == io_wptr_0 ? io_dataIn_0 : table_19; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_288 = 5'h14 == io_wptr_0 ? io_dataIn_0 : table_20; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_289 = 5'h15 == io_wptr_0 ? io_dataIn_0 : table_21; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_290 = 5'h16 == io_wptr_0 ? io_dataIn_0 : table_22; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_291 = 5'h17 == io_wptr_0 ? io_dataIn_0 : table_23; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_292 = 5'h18 == io_wptr_0 ? io_dataIn_0 : table_24; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_293 = 5'h19 == io_wptr_0 ? io_dataIn_0 : table_25; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_294 = 5'h1a == io_wptr_0 ? io_dataIn_0 : table_26; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_295 = 5'h1b == io_wptr_0 ? io_dataIn_0 : table_27; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_296 = 5'h1c == io_wptr_0 ? io_dataIn_0 : table_28; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_297 = 5'h1d == io_wptr_0 ? io_dataIn_0 : table_29; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_298 = 5'h1e == io_wptr_0 ? io_dataIn_0 : table_30; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_299 = 5'h1f == io_wptr_0 ? io_dataIn_0 : table_31; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_300 = 5'h0 == io_wptr_1 ? io_dataIn_1 : _GEN_268; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_301 = 5'h1 == io_wptr_1 ? io_dataIn_1 : _GEN_269; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_302 = 5'h2 == io_wptr_1 ? io_dataIn_1 : _GEN_270; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_303 = 5'h3 == io_wptr_1 ? io_dataIn_1 : _GEN_271; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_304 = 5'h4 == io_wptr_1 ? io_dataIn_1 : _GEN_272; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_305 = 5'h5 == io_wptr_1 ? io_dataIn_1 : _GEN_273; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_306 = 5'h6 == io_wptr_1 ? io_dataIn_1 : _GEN_274; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_307 = 5'h7 == io_wptr_1 ? io_dataIn_1 : _GEN_275; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_308 = 5'h8 == io_wptr_1 ? io_dataIn_1 : _GEN_276; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_309 = 5'h9 == io_wptr_1 ? io_dataIn_1 : _GEN_277; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_310 = 5'ha == io_wptr_1 ? io_dataIn_1 : _GEN_278; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_311 = 5'hb == io_wptr_1 ? io_dataIn_1 : _GEN_279; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_312 = 5'hc == io_wptr_1 ? io_dataIn_1 : _GEN_280; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_313 = 5'hd == io_wptr_1 ? io_dataIn_1 : _GEN_281; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_314 = 5'he == io_wptr_1 ? io_dataIn_1 : _GEN_282; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_315 = 5'hf == io_wptr_1 ? io_dataIn_1 : _GEN_283; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_316 = 5'h10 == io_wptr_1 ? io_dataIn_1 : _GEN_284; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_317 = 5'h11 == io_wptr_1 ? io_dataIn_1 : _GEN_285; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_318 = 5'h12 == io_wptr_1 ? io_dataIn_1 : _GEN_286; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_319 = 5'h13 == io_wptr_1 ? io_dataIn_1 : _GEN_287; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_320 = 5'h14 == io_wptr_1 ? io_dataIn_1 : _GEN_288; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_321 = 5'h15 == io_wptr_1 ? io_dataIn_1 : _GEN_289; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_322 = 5'h16 == io_wptr_1 ? io_dataIn_1 : _GEN_290; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_323 = 5'h17 == io_wptr_1 ? io_dataIn_1 : _GEN_291; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_324 = 5'h18 == io_wptr_1 ? io_dataIn_1 : _GEN_292; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_325 = 5'h19 == io_wptr_1 ? io_dataIn_1 : _GEN_293; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_326 = 5'h1a == io_wptr_1 ? io_dataIn_1 : _GEN_294; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_327 = 5'h1b == io_wptr_1 ? io_dataIn_1 : _GEN_295; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_328 = 5'h1c == io_wptr_1 ? io_dataIn_1 : _GEN_296; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_329 = 5'h1d == io_wptr_1 ? io_dataIn_1 : _GEN_297; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_330 = 5'h1e == io_wptr_1 ? io_dataIn_1 : _GEN_298; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_331 = 5'h1f == io_wptr_1 ? io_dataIn_1 : _GEN_299; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_364 = 5'h0 == io_wptr_1 ? io_dataIn_1 : table_0; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_365 = 5'h1 == io_wptr_1 ? io_dataIn_1 : table_1; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_366 = 5'h2 == io_wptr_1 ? io_dataIn_1 : table_2; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_367 = 5'h3 == io_wptr_1 ? io_dataIn_1 : table_3; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_368 = 5'h4 == io_wptr_1 ? io_dataIn_1 : table_4; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_369 = 5'h5 == io_wptr_1 ? io_dataIn_1 : table_5; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_370 = 5'h6 == io_wptr_1 ? io_dataIn_1 : table_6; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_371 = 5'h7 == io_wptr_1 ? io_dataIn_1 : table_7; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_372 = 5'h8 == io_wptr_1 ? io_dataIn_1 : table_8; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_373 = 5'h9 == io_wptr_1 ? io_dataIn_1 : table_9; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_374 = 5'ha == io_wptr_1 ? io_dataIn_1 : table_10; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_375 = 5'hb == io_wptr_1 ? io_dataIn_1 : table_11; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_376 = 5'hc == io_wptr_1 ? io_dataIn_1 : table_12; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_377 = 5'hd == io_wptr_1 ? io_dataIn_1 : table_13; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_378 = 5'he == io_wptr_1 ? io_dataIn_1 : table_14; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_379 = 5'hf == io_wptr_1 ? io_dataIn_1 : table_15; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_380 = 5'h10 == io_wptr_1 ? io_dataIn_1 : table_16; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_381 = 5'h11 == io_wptr_1 ? io_dataIn_1 : table_17; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_382 = 5'h12 == io_wptr_1 ? io_dataIn_1 : table_18; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_383 = 5'h13 == io_wptr_1 ? io_dataIn_1 : table_19; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_384 = 5'h14 == io_wptr_1 ? io_dataIn_1 : table_20; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_385 = 5'h15 == io_wptr_1 ? io_dataIn_1 : table_21; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_386 = 5'h16 == io_wptr_1 ? io_dataIn_1 : table_22; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_387 = 5'h17 == io_wptr_1 ? io_dataIn_1 : table_23; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_388 = 5'h18 == io_wptr_1 ? io_dataIn_1 : table_24; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_389 = 5'h19 == io_wptr_1 ? io_dataIn_1 : table_25; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_390 = 5'h1a == io_wptr_1 ? io_dataIn_1 : table_26; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_391 = 5'h1b == io_wptr_1 ? io_dataIn_1 : table_27; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_392 = 5'h1c == io_wptr_1 ? io_dataIn_1 : table_28; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_393 = 5'h1d == io_wptr_1 ? io_dataIn_1 : table_29; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_394 = 5'h1e == io_wptr_1 ? io_dataIn_1 : table_30; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_395 = 5'h1f == io_wptr_1 ? io_dataIn_1 : table_31; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_396 = io_writeFlag_1 ? _GEN_364 : table_0; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_397 = io_writeFlag_1 ? _GEN_365 : table_1; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_398 = io_writeFlag_1 ? _GEN_366 : table_2; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_399 = io_writeFlag_1 ? _GEN_367 : table_3; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_400 = io_writeFlag_1 ? _GEN_368 : table_4; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_401 = io_writeFlag_1 ? _GEN_369 : table_5; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_402 = io_writeFlag_1 ? _GEN_370 : table_6; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_403 = io_writeFlag_1 ? _GEN_371 : table_7; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_404 = io_writeFlag_1 ? _GEN_372 : table_8; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_405 = io_writeFlag_1 ? _GEN_373 : table_9; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_406 = io_writeFlag_1 ? _GEN_374 : table_10; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_407 = io_writeFlag_1 ? _GEN_375 : table_11; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_408 = io_writeFlag_1 ? _GEN_376 : table_12; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_409 = io_writeFlag_1 ? _GEN_377 : table_13; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_410 = io_writeFlag_1 ? _GEN_378 : table_14; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_411 = io_writeFlag_1 ? _GEN_379 : table_15; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_412 = io_writeFlag_1 ? _GEN_380 : table_16; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_413 = io_writeFlag_1 ? _GEN_381 : table_17; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_414 = io_writeFlag_1 ? _GEN_382 : table_18; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_415 = io_writeFlag_1 ? _GEN_383 : table_19; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_416 = io_writeFlag_1 ? _GEN_384 : table_20; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_417 = io_writeFlag_1 ? _GEN_385 : table_21; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_418 = io_writeFlag_1 ? _GEN_386 : table_22; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_419 = io_writeFlag_1 ? _GEN_387 : table_23; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_420 = io_writeFlag_1 ? _GEN_388 : table_24; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_421 = io_writeFlag_1 ? _GEN_389 : table_25; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_422 = io_writeFlag_1 ? _GEN_390 : table_26; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_423 = io_writeFlag_1 ? _GEN_391 : table_27; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_424 = io_writeFlag_1 ? _GEN_392 : table_28; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_425 = io_writeFlag_1 ? _GEN_393 : table_29; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_426 = io_writeFlag_1 ? _GEN_394 : table_30; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_427 = io_writeFlag_1 ? _GEN_395 : table_31; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_428 = io_writeFlag_0 ? _GEN_268 : _GEN_396; // @[util.scala 85:30]
  wire [31:0] _GEN_429 = io_writeFlag_0 ? _GEN_269 : _GEN_397; // @[util.scala 85:30]
  wire [31:0] _GEN_430 = io_writeFlag_0 ? _GEN_270 : _GEN_398; // @[util.scala 85:30]
  wire [31:0] _GEN_431 = io_writeFlag_0 ? _GEN_271 : _GEN_399; // @[util.scala 85:30]
  wire [31:0] _GEN_432 = io_writeFlag_0 ? _GEN_272 : _GEN_400; // @[util.scala 85:30]
  wire [31:0] _GEN_433 = io_writeFlag_0 ? _GEN_273 : _GEN_401; // @[util.scala 85:30]
  wire [31:0] _GEN_434 = io_writeFlag_0 ? _GEN_274 : _GEN_402; // @[util.scala 85:30]
  wire [31:0] _GEN_435 = io_writeFlag_0 ? _GEN_275 : _GEN_403; // @[util.scala 85:30]
  wire [31:0] _GEN_436 = io_writeFlag_0 ? _GEN_276 : _GEN_404; // @[util.scala 85:30]
  wire [31:0] _GEN_437 = io_writeFlag_0 ? _GEN_277 : _GEN_405; // @[util.scala 85:30]
  wire [31:0] _GEN_438 = io_writeFlag_0 ? _GEN_278 : _GEN_406; // @[util.scala 85:30]
  wire [31:0] _GEN_439 = io_writeFlag_0 ? _GEN_279 : _GEN_407; // @[util.scala 85:30]
  wire [31:0] _GEN_440 = io_writeFlag_0 ? _GEN_280 : _GEN_408; // @[util.scala 85:30]
  wire [31:0] _GEN_441 = io_writeFlag_0 ? _GEN_281 : _GEN_409; // @[util.scala 85:30]
  wire [31:0] _GEN_442 = io_writeFlag_0 ? _GEN_282 : _GEN_410; // @[util.scala 85:30]
  wire [31:0] _GEN_443 = io_writeFlag_0 ? _GEN_283 : _GEN_411; // @[util.scala 85:30]
  wire [31:0] _GEN_444 = io_writeFlag_0 ? _GEN_284 : _GEN_412; // @[util.scala 85:30]
  wire [31:0] _GEN_445 = io_writeFlag_0 ? _GEN_285 : _GEN_413; // @[util.scala 85:30]
  wire [31:0] _GEN_446 = io_writeFlag_0 ? _GEN_286 : _GEN_414; // @[util.scala 85:30]
  wire [31:0] _GEN_447 = io_writeFlag_0 ? _GEN_287 : _GEN_415; // @[util.scala 85:30]
  wire [31:0] _GEN_448 = io_writeFlag_0 ? _GEN_288 : _GEN_416; // @[util.scala 85:30]
  wire [31:0] _GEN_449 = io_writeFlag_0 ? _GEN_289 : _GEN_417; // @[util.scala 85:30]
  wire [31:0] _GEN_450 = io_writeFlag_0 ? _GEN_290 : _GEN_418; // @[util.scala 85:30]
  wire [31:0] _GEN_451 = io_writeFlag_0 ? _GEN_291 : _GEN_419; // @[util.scala 85:30]
  wire [31:0] _GEN_452 = io_writeFlag_0 ? _GEN_292 : _GEN_420; // @[util.scala 85:30]
  wire [31:0] _GEN_453 = io_writeFlag_0 ? _GEN_293 : _GEN_421; // @[util.scala 85:30]
  wire [31:0] _GEN_454 = io_writeFlag_0 ? _GEN_294 : _GEN_422; // @[util.scala 85:30]
  wire [31:0] _GEN_455 = io_writeFlag_0 ? _GEN_295 : _GEN_423; // @[util.scala 85:30]
  wire [31:0] _GEN_456 = io_writeFlag_0 ? _GEN_296 : _GEN_424; // @[util.scala 85:30]
  wire [31:0] _GEN_457 = io_writeFlag_0 ? _GEN_297 : _GEN_425; // @[util.scala 85:30]
  wire [31:0] _GEN_458 = io_writeFlag_0 ? _GEN_298 : _GEN_426; // @[util.scala 85:30]
  wire [31:0] _GEN_459 = io_writeFlag_0 ? _GEN_299 : _GEN_427; // @[util.scala 85:30]
  wire [31:0] _GEN_460 = _T_7 ? _GEN_300 : _GEN_428; // @[util.scala 82:39]
  wire [31:0] _GEN_461 = _T_7 ? _GEN_301 : _GEN_429; // @[util.scala 82:39]
  wire [31:0] _GEN_462 = _T_7 ? _GEN_302 : _GEN_430; // @[util.scala 82:39]
  wire [31:0] _GEN_463 = _T_7 ? _GEN_303 : _GEN_431; // @[util.scala 82:39]
  wire [31:0] _GEN_464 = _T_7 ? _GEN_304 : _GEN_432; // @[util.scala 82:39]
  wire [31:0] _GEN_465 = _T_7 ? _GEN_305 : _GEN_433; // @[util.scala 82:39]
  wire [31:0] _GEN_466 = _T_7 ? _GEN_306 : _GEN_434; // @[util.scala 82:39]
  wire [31:0] _GEN_467 = _T_7 ? _GEN_307 : _GEN_435; // @[util.scala 82:39]
  wire [31:0] _GEN_468 = _T_7 ? _GEN_308 : _GEN_436; // @[util.scala 82:39]
  wire [31:0] _GEN_469 = _T_7 ? _GEN_309 : _GEN_437; // @[util.scala 82:39]
  wire [31:0] _GEN_470 = _T_7 ? _GEN_310 : _GEN_438; // @[util.scala 82:39]
  wire [31:0] _GEN_471 = _T_7 ? _GEN_311 : _GEN_439; // @[util.scala 82:39]
  wire [31:0] _GEN_472 = _T_7 ? _GEN_312 : _GEN_440; // @[util.scala 82:39]
  wire [31:0] _GEN_473 = _T_7 ? _GEN_313 : _GEN_441; // @[util.scala 82:39]
  wire [31:0] _GEN_474 = _T_7 ? _GEN_314 : _GEN_442; // @[util.scala 82:39]
  wire [31:0] _GEN_475 = _T_7 ? _GEN_315 : _GEN_443; // @[util.scala 82:39]
  wire [31:0] _GEN_476 = _T_7 ? _GEN_316 : _GEN_444; // @[util.scala 82:39]
  wire [31:0] _GEN_477 = _T_7 ? _GEN_317 : _GEN_445; // @[util.scala 82:39]
  wire [31:0] _GEN_478 = _T_7 ? _GEN_318 : _GEN_446; // @[util.scala 82:39]
  wire [31:0] _GEN_479 = _T_7 ? _GEN_319 : _GEN_447; // @[util.scala 82:39]
  wire [31:0] _GEN_480 = _T_7 ? _GEN_320 : _GEN_448; // @[util.scala 82:39]
  wire [31:0] _GEN_481 = _T_7 ? _GEN_321 : _GEN_449; // @[util.scala 82:39]
  wire [31:0] _GEN_482 = _T_7 ? _GEN_322 : _GEN_450; // @[util.scala 82:39]
  wire [31:0] _GEN_483 = _T_7 ? _GEN_323 : _GEN_451; // @[util.scala 82:39]
  wire [31:0] _GEN_484 = _T_7 ? _GEN_324 : _GEN_452; // @[util.scala 82:39]
  wire [31:0] _GEN_485 = _T_7 ? _GEN_325 : _GEN_453; // @[util.scala 82:39]
  wire [31:0] _GEN_486 = _T_7 ? _GEN_326 : _GEN_454; // @[util.scala 82:39]
  wire [31:0] _GEN_487 = _T_7 ? _GEN_327 : _GEN_455; // @[util.scala 82:39]
  wire [31:0] _GEN_488 = _T_7 ? _GEN_328 : _GEN_456; // @[util.scala 82:39]
  wire [31:0] _GEN_489 = _T_7 ? _GEN_329 : _GEN_457; // @[util.scala 82:39]
  wire [31:0] _GEN_490 = _T_7 ? _GEN_330 : _GEN_458; // @[util.scala 82:39]
  wire [31:0] _GEN_491 = _T_7 ? _GEN_331 : _GEN_459; // @[util.scala 82:39]
  wire [31:0] _GEN_492 = wvalid ? _GEN_12 : _GEN_460; // @[util.scala 80:21]
  wire [31:0] _GEN_493 = wvalid ? _GEN_13 : _GEN_461; // @[util.scala 80:21]
  wire [31:0] _GEN_494 = wvalid ? _GEN_14 : _GEN_462; // @[util.scala 80:21]
  wire [31:0] _GEN_495 = wvalid ? _GEN_15 : _GEN_463; // @[util.scala 80:21]
  wire [31:0] _GEN_496 = wvalid ? _GEN_16 : _GEN_464; // @[util.scala 80:21]
  wire [31:0] _GEN_497 = wvalid ? _GEN_17 : _GEN_465; // @[util.scala 80:21]
  wire [31:0] _GEN_498 = wvalid ? _GEN_18 : _GEN_466; // @[util.scala 80:21]
  wire [31:0] _GEN_499 = wvalid ? _GEN_19 : _GEN_467; // @[util.scala 80:21]
  wire [31:0] _GEN_500 = wvalid ? _GEN_20 : _GEN_468; // @[util.scala 80:21]
  wire [31:0] _GEN_501 = wvalid ? _GEN_21 : _GEN_469; // @[util.scala 80:21]
  wire [31:0] _GEN_502 = wvalid ? _GEN_22 : _GEN_470; // @[util.scala 80:21]
  wire [31:0] _GEN_503 = wvalid ? _GEN_23 : _GEN_471; // @[util.scala 80:21]
  wire [31:0] _GEN_504 = wvalid ? _GEN_24 : _GEN_472; // @[util.scala 80:21]
  wire [31:0] _GEN_505 = wvalid ? _GEN_25 : _GEN_473; // @[util.scala 80:21]
  wire [31:0] _GEN_506 = wvalid ? _GEN_26 : _GEN_474; // @[util.scala 80:21]
  wire [31:0] _GEN_507 = wvalid ? _GEN_27 : _GEN_475; // @[util.scala 80:21]
  wire [31:0] _GEN_508 = wvalid ? _GEN_28 : _GEN_476; // @[util.scala 80:21]
  wire [31:0] _GEN_509 = wvalid ? _GEN_29 : _GEN_477; // @[util.scala 80:21]
  wire [31:0] _GEN_510 = wvalid ? _GEN_30 : _GEN_478; // @[util.scala 80:21]
  wire [31:0] _GEN_511 = wvalid ? _GEN_31 : _GEN_479; // @[util.scala 80:21]
  wire [31:0] _GEN_512 = wvalid ? _GEN_32 : _GEN_480; // @[util.scala 80:21]
  wire [31:0] _GEN_513 = wvalid ? _GEN_33 : _GEN_481; // @[util.scala 80:21]
  wire [31:0] _GEN_514 = wvalid ? _GEN_34 : _GEN_482; // @[util.scala 80:21]
  wire [31:0] _GEN_515 = wvalid ? _GEN_35 : _GEN_483; // @[util.scala 80:21]
  wire [31:0] _GEN_516 = wvalid ? _GEN_36 : _GEN_484; // @[util.scala 80:21]
  wire [31:0] _GEN_517 = wvalid ? _GEN_37 : _GEN_485; // @[util.scala 80:21]
  wire [31:0] _GEN_518 = wvalid ? _GEN_38 : _GEN_486; // @[util.scala 80:21]
  wire [31:0] _GEN_519 = wvalid ? _GEN_39 : _GEN_487; // @[util.scala 80:21]
  wire [31:0] _GEN_520 = wvalid ? _GEN_40 : _GEN_488; // @[util.scala 80:21]
  wire [31:0] _GEN_521 = wvalid ? _GEN_41 : _GEN_489; // @[util.scala 80:21]
  wire [31:0] _GEN_522 = wvalid ? _GEN_42 : _GEN_490; // @[util.scala 80:21]
  wire [31:0] _GEN_523 = wvalid ? _GEN_43 : _GEN_491; // @[util.scala 80:21]
  reg [4:0] eraddr; // @[util.scala 92:19]
  wire [31:0] _GEN_622 = 5'h1 == eraddr ? table_1 : table_0; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_623 = 5'h2 == eraddr ? table_2 : _GEN_622; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_624 = 5'h3 == eraddr ? table_3 : _GEN_623; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_625 = 5'h4 == eraddr ? table_4 : _GEN_624; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_626 = 5'h5 == eraddr ? table_5 : _GEN_625; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_627 = 5'h6 == eraddr ? table_6 : _GEN_626; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_628 = 5'h7 == eraddr ? table_7 : _GEN_627; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_629 = 5'h8 == eraddr ? table_8 : _GEN_628; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_630 = 5'h9 == eraddr ? table_9 : _GEN_629; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_631 = 5'ha == eraddr ? table_10 : _GEN_630; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_632 = 5'hb == eraddr ? table_11 : _GEN_631; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_633 = 5'hc == eraddr ? table_12 : _GEN_632; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_634 = 5'hd == eraddr ? table_13 : _GEN_633; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_635 = 5'he == eraddr ? table_14 : _GEN_634; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_636 = 5'hf == eraddr ? table_15 : _GEN_635; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_637 = 5'h10 == eraddr ? table_16 : _GEN_636; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_638 = 5'h11 == eraddr ? table_17 : _GEN_637; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_639 = 5'h12 == eraddr ? table_18 : _GEN_638; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_640 = 5'h13 == eraddr ? table_19 : _GEN_639; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_641 = 5'h14 == eraddr ? table_20 : _GEN_640; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_642 = 5'h15 == eraddr ? table_21 : _GEN_641; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_643 = 5'h16 == eraddr ? table_22 : _GEN_642; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_644 = 5'h17 == eraddr ? table_23 : _GEN_643; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_645 = 5'h18 == eraddr ? table_24 : _GEN_644; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_646 = 5'h19 == eraddr ? table_25 : _GEN_645; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_647 = 5'h1a == eraddr ? table_26 : _GEN_646; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_648 = 5'h1b == eraddr ? table_27 : _GEN_647; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_649 = 5'h1c == eraddr ? table_28 : _GEN_648; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_650 = 5'h1d == eraddr ? table_29 : _GEN_649; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_651 = 5'h1e == eraddr ? table_30 : _GEN_650; // @[util.scala 99:16 util.scala 99:16]
  assign io_data_0 = table_0; // @[util.scala 53:11]
  assign io_data_1 = table_1; // @[util.scala 53:11]
  assign io_data_2 = table_2; // @[util.scala 53:11]
  assign io_data_3 = table_3; // @[util.scala 53:11]
  assign io_data_4 = table_4; // @[util.scala 53:11]
  assign io_data_7 = table_7; // @[util.scala 53:11]
  assign io_data_12 = table_12; // @[util.scala 53:11]
  assign io_data_13 = table_13; // @[util.scala 53:11]
  assign io_data_16 = table_16; // @[util.scala 53:11]
  assign io_data_17 = table_17; // @[util.scala 53:11]
  assign io_data_18 = table_18; // @[util.scala 53:11]
  assign io_data_19 = table_19; // @[util.scala 53:11]
  assign io_data_20 = table_20; // @[util.scala 53:11]
  assign io_data_21 = table_21; // @[util.scala 53:11]
  assign io_data_22 = table_22; // @[util.scala 53:11]
  assign io_data_23 = table_23; // @[util.scala 53:11]
  assign io_data_24 = table_24; // @[util.scala 53:11]
  assign io_data_25 = table_25; // @[util.scala 53:11]
  assign io_data_26 = table_26; // @[util.scala 53:11]
  assign io_data_27 = table_27; // @[util.scala 53:11]
  assign io_data_28 = table_28; // @[util.scala 53:11]
  assign io_data_29 = table_29; // @[util.scala 53:11]
  assign config_awready = status == 3'h0; // @[util.scala 55:28]
  assign config_arready = status == 3'h0; // @[util.scala 56:28]
  assign config_wready = status == 3'h1; // @[util.scala 54:27]
  assign config_rdata = 5'h1f == eraddr ? table_31 : _GEN_651; // @[util.scala 99:16 util.scala 99:16]
  assign config_rvalid = status == 3'h5; // @[util.scala 57:27]
  assign config_bvalid = status == 3'h3; // @[util.scala 58:27]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 16:22]
      table_0 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h0 == io_wptr_1) begin // @[util.scala 73:23]
        table_0 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_0 <= _GEN_44;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_0 <= _GEN_44;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_0 <= _GEN_204;
    end else begin
      table_0 <= _GEN_492;
    end
    if (reset) begin // @[util.scala 16:22]
      table_1 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1 == io_wptr_1) begin // @[util.scala 73:23]
        table_1 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_1 <= _GEN_45;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_1 <= _GEN_45;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_1 <= _GEN_205;
    end else begin
      table_1 <= _GEN_493;
    end
    if (reset) begin // @[util.scala 16:22]
      table_2 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h2 == io_wptr_1) begin // @[util.scala 73:23]
        table_2 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_2 <= _GEN_46;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_2 <= _GEN_46;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_2 <= _GEN_206;
    end else begin
      table_2 <= _GEN_494;
    end
    if (reset) begin // @[util.scala 16:22]
      table_3 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h3 == io_wptr_1) begin // @[util.scala 73:23]
        table_3 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_3 <= _GEN_47;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_3 <= _GEN_47;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_3 <= _GEN_207;
    end else begin
      table_3 <= _GEN_495;
    end
    if (reset) begin // @[util.scala 16:22]
      table_4 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h4 == io_wptr_1) begin // @[util.scala 73:23]
        table_4 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_4 <= _GEN_48;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_4 <= _GEN_48;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_4 <= _GEN_208;
    end else begin
      table_4 <= _GEN_496;
    end
    if (reset) begin // @[util.scala 16:22]
      table_5 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h5 == io_wptr_1) begin // @[util.scala 73:23]
        table_5 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_5 <= _GEN_49;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_5 <= _GEN_49;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_5 <= _GEN_209;
    end else begin
      table_5 <= _GEN_497;
    end
    if (reset) begin // @[util.scala 16:22]
      table_6 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h6 == io_wptr_1) begin // @[util.scala 73:23]
        table_6 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_6 <= _GEN_50;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_6 <= _GEN_50;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_6 <= _GEN_210;
    end else begin
      table_6 <= _GEN_498;
    end
    if (reset) begin // @[util.scala 16:22]
      table_7 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h7 == io_wptr_1) begin // @[util.scala 73:23]
        table_7 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_7 <= _GEN_51;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_7 <= _GEN_51;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_7 <= _GEN_211;
    end else begin
      table_7 <= _GEN_499;
    end
    if (reset) begin // @[util.scala 16:22]
      table_8 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h8 == io_wptr_1) begin // @[util.scala 73:23]
        table_8 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_8 <= _GEN_52;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_8 <= _GEN_52;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_8 <= _GEN_212;
    end else begin
      table_8 <= _GEN_500;
    end
    if (reset) begin // @[util.scala 16:22]
      table_9 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h9 == io_wptr_1) begin // @[util.scala 73:23]
        table_9 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_9 <= _GEN_53;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_9 <= _GEN_53;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_9 <= _GEN_213;
    end else begin
      table_9 <= _GEN_501;
    end
    if (reset) begin // @[util.scala 16:22]
      table_10 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'ha == io_wptr_1) begin // @[util.scala 73:23]
        table_10 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_10 <= _GEN_54;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_10 <= _GEN_54;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_10 <= _GEN_214;
    end else begin
      table_10 <= _GEN_502;
    end
    if (reset) begin // @[util.scala 16:22]
      table_11 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hb == io_wptr_1) begin // @[util.scala 73:23]
        table_11 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_11 <= _GEN_55;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_11 <= _GEN_55;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_11 <= _GEN_215;
    end else begin
      table_11 <= _GEN_503;
    end
    if (reset) begin // @[util.scala 16:22]
      table_12 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hc == io_wptr_1) begin // @[util.scala 73:23]
        table_12 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_12 <= _GEN_56;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_12 <= _GEN_56;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_12 <= _GEN_216;
    end else begin
      table_12 <= _GEN_504;
    end
    if (reset) begin // @[util.scala 16:22]
      table_13 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hd == io_wptr_1) begin // @[util.scala 73:23]
        table_13 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_13 <= _GEN_57;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_13 <= _GEN_57;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_13 <= _GEN_217;
    end else begin
      table_13 <= _GEN_505;
    end
    if (reset) begin // @[util.scala 16:22]
      table_14 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'he == io_wptr_1) begin // @[util.scala 73:23]
        table_14 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_14 <= _GEN_58;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_14 <= _GEN_58;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_14 <= _GEN_218;
    end else begin
      table_14 <= _GEN_506;
    end
    if (reset) begin // @[util.scala 16:22]
      table_15 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hf == io_wptr_1) begin // @[util.scala 73:23]
        table_15 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_15 <= _GEN_59;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_15 <= _GEN_59;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_15 <= _GEN_219;
    end else begin
      table_15 <= _GEN_507;
    end
    if (reset) begin // @[util.scala 16:22]
      table_16 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h10 == io_wptr_1) begin // @[util.scala 73:23]
        table_16 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_16 <= _GEN_60;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_16 <= _GEN_60;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_16 <= _GEN_220;
    end else begin
      table_16 <= _GEN_508;
    end
    if (reset) begin // @[util.scala 16:22]
      table_17 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h11 == io_wptr_1) begin // @[util.scala 73:23]
        table_17 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_17 <= _GEN_61;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_17 <= _GEN_61;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_17 <= _GEN_221;
    end else begin
      table_17 <= _GEN_509;
    end
    if (reset) begin // @[util.scala 16:22]
      table_18 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h12 == io_wptr_1) begin // @[util.scala 73:23]
        table_18 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_18 <= _GEN_62;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_18 <= _GEN_62;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_18 <= _GEN_222;
    end else begin
      table_18 <= _GEN_510;
    end
    if (reset) begin // @[util.scala 16:22]
      table_19 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h13 == io_wptr_1) begin // @[util.scala 73:23]
        table_19 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_19 <= _GEN_63;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_19 <= _GEN_63;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_19 <= _GEN_223;
    end else begin
      table_19 <= _GEN_511;
    end
    if (reset) begin // @[util.scala 16:22]
      table_20 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h14 == io_wptr_1) begin // @[util.scala 73:23]
        table_20 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_20 <= _GEN_64;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_20 <= _GEN_64;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_20 <= _GEN_224;
    end else begin
      table_20 <= _GEN_512;
    end
    if (reset) begin // @[util.scala 16:22]
      table_21 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h15 == io_wptr_1) begin // @[util.scala 73:23]
        table_21 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_21 <= _GEN_65;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_21 <= _GEN_65;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_21 <= _GEN_225;
    end else begin
      table_21 <= _GEN_513;
    end
    if (reset) begin // @[util.scala 16:22]
      table_22 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h16 == io_wptr_1) begin // @[util.scala 73:23]
        table_22 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_22 <= _GEN_66;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_22 <= _GEN_66;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_22 <= _GEN_226;
    end else begin
      table_22 <= _GEN_514;
    end
    if (reset) begin // @[util.scala 16:22]
      table_23 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h17 == io_wptr_1) begin // @[util.scala 73:23]
        table_23 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_23 <= _GEN_67;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_23 <= _GEN_67;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_23 <= _GEN_227;
    end else begin
      table_23 <= _GEN_515;
    end
    if (reset) begin // @[util.scala 16:22]
      table_24 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h18 == io_wptr_1) begin // @[util.scala 73:23]
        table_24 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_24 <= _GEN_68;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_24 <= _GEN_68;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_24 <= _GEN_228;
    end else begin
      table_24 <= _GEN_516;
    end
    if (reset) begin // @[util.scala 16:22]
      table_25 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h19 == io_wptr_1) begin // @[util.scala 73:23]
        table_25 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_25 <= _GEN_69;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_25 <= _GEN_69;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_25 <= _GEN_229;
    end else begin
      table_25 <= _GEN_517;
    end
    if (reset) begin // @[util.scala 16:22]
      table_26 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1a == io_wptr_1) begin // @[util.scala 73:23]
        table_26 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_26 <= _GEN_70;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_26 <= _GEN_70;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_26 <= _GEN_230;
    end else begin
      table_26 <= _GEN_518;
    end
    if (reset) begin // @[util.scala 16:22]
      table_27 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1b == io_wptr_1) begin // @[util.scala 73:23]
        table_27 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_27 <= _GEN_71;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_27 <= _GEN_71;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_27 <= _GEN_231;
    end else begin
      table_27 <= _GEN_519;
    end
    if (reset) begin // @[util.scala 16:22]
      table_28 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1c == io_wptr_1) begin // @[util.scala 73:23]
        table_28 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_28 <= _GEN_72;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_28 <= _GEN_72;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_28 <= _GEN_232;
    end else begin
      table_28 <= _GEN_520;
    end
    if (reset) begin // @[util.scala 16:22]
      table_29 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1d == io_wptr_1) begin // @[util.scala 73:23]
        table_29 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_29 <= _GEN_73;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_29 <= _GEN_73;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_29 <= _GEN_233;
    end else begin
      table_29 <= _GEN_521;
    end
    if (reset) begin // @[util.scala 16:22]
      table_30 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1e == io_wptr_1) begin // @[util.scala 73:23]
        table_30 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_30 <= _GEN_74;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_30 <= _GEN_74;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_30 <= _GEN_234;
    end else begin
      table_30 <= _GEN_522;
    end
    if (reset) begin // @[util.scala 16:22]
      table_31 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1f == io_wptr_1) begin // @[util.scala 73:23]
        table_31 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_31 <= _GEN_75;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_31 <= _GEN_75;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_31 <= _GEN_235;
    end else begin
      table_31 <= _GEN_523;
    end
    if (reset) begin // @[util.scala 26:23]
      status <= 3'h0; // @[util.scala 26:23]
    end else if (status == 3'h0) begin // @[util.scala 28:28]
      if (config_awvalid) begin // @[util.scala 29:25]
        status <= 3'h1; // @[util.scala 30:14]
      end else if (config_arvalid) begin // @[util.scala 31:31]
        status <= 3'h4; // @[util.scala 32:14]
      end
    end else if (status == 3'h1) begin // @[util.scala 34:35]
      if (config_wvalid) begin // @[util.scala 35:24]
        status <= 3'h2; // @[util.scala 36:14]
      end
    end else if (status == 3'h2) begin // @[util.scala 38:34]
      status <= 3'h3; // @[util.scala 39:12]
    end else begin
      status <= _GEN_7;
    end
    if (config_awvalid & config_awready) begin // @[util.scala 66:41]
      ewaddr <= config_awaddr[6:2]; // @[util.scala 67:12]
    end
    if (config_arvalid & config_arready) begin // @[util.scala 93:41]
      eraddr <= config_araddr[6:2]; // @[util.scala 94:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  table_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  table_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  table_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  table_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  table_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  table_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  table_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  table_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  table_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  table_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  table_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  table_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  table_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  table_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  table_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  table_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  table_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  table_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  table_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  table_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  table_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  table_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  table_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  table_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  table_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  table_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  table_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  table_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  table_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  table_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  table_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  table_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  status = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  ewaddr = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  eraddr = _RAND_34[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module controller(
  input         clock,
  input         reset,
  output [31:0] io_data_0,
  output [31:0] io_data_1,
  output [31:0] io_data_2,
  output [31:0] io_data_3,
  output [31:0] io_data_4,
  output [31:0] io_data_7,
  output [31:0] io_data_16,
  output [31:0] io_data_17,
  output [31:0] io_data_18,
  output [31:0] io_data_19,
  output [31:0] io_data_20,
  output [31:0] io_data_21,
  output [31:0] io_data_22,
  output [31:0] io_data_23,
  output [31:0] io_data_24,
  output [31:0] io_data_25,
  output [31:0] io_data_26,
  output [31:0] io_data_27,
  output [31:0] io_data_28,
  output [31:0] io_data_29,
  input         io_fin_0,
  input         io_fin_1,
  input         io_fin_2,
  input         io_fin_3,
  input         io_fin_4,
  input         io_fin_5,
  input         io_fin_6,
  input         io_fin_7,
  input         io_fin_8,
  input         io_fin_9,
  input         io_fin_10,
  input         io_fin_11,
  input         io_fin_12,
  input         io_fin_13,
  input         io_fin_14,
  input         io_fin_15,
  input         io_fin_16,
  input         io_fin_17,
  input         io_fin_18,
  input         io_fin_19,
  output        io_signal,
  output        io_start,
  output [31:0] io_level,
  input  [63:0] io_traveled_edges,
  input  [63:0] io_config_awaddr,
  input         io_config_awvalid,
  output        io_config_awready,
  input  [63:0] io_config_araddr,
  input         io_config_arvalid,
  output        io_config_arready,
  input  [31:0] io_config_wdata,
  input         io_config_wvalid,
  output        io_config_wready,
  output [31:0] io_config_rdata,
  output        io_config_rvalid,
  input         io_config_rready,
  output        io_config_bvalid,
  input         io_config_bready,
  output        io_flush_cache,
  input         io_flush_cache_end,
  input         io_signal_ack
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  wire  controls_clock; // @[BFS.scala 1125:24]
  wire  controls_reset; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_0; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_1; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_2; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_3; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_4; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_7; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_12; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_13; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_16; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_17; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_18; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_19; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_20; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_21; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_22; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_23; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_24; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_25; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_26; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_27; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_28; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_data_29; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_dataIn_0; // @[BFS.scala 1125:24]
  wire [31:0] controls_io_dataIn_1; // @[BFS.scala 1125:24]
  wire  controls_io_writeFlag_0; // @[BFS.scala 1125:24]
  wire  controls_io_writeFlag_1; // @[BFS.scala 1125:24]
  wire [4:0] controls_io_wptr_0; // @[BFS.scala 1125:24]
  wire [4:0] controls_io_wptr_1; // @[BFS.scala 1125:24]
  wire [63:0] controls_config_awaddr; // @[BFS.scala 1125:24]
  wire  controls_config_awvalid; // @[BFS.scala 1125:24]
  wire  controls_config_awready; // @[BFS.scala 1125:24]
  wire [63:0] controls_config_araddr; // @[BFS.scala 1125:24]
  wire  controls_config_arvalid; // @[BFS.scala 1125:24]
  wire  controls_config_arready; // @[BFS.scala 1125:24]
  wire [31:0] controls_config_wdata; // @[BFS.scala 1125:24]
  wire  controls_config_wvalid; // @[BFS.scala 1125:24]
  wire  controls_config_wready; // @[BFS.scala 1125:24]
  wire [31:0] controls_config_rdata; // @[BFS.scala 1125:24]
  wire  controls_config_rvalid; // @[BFS.scala 1125:24]
  wire  controls_config_rready; // @[BFS.scala 1125:24]
  wire  controls_config_bvalid; // @[BFS.scala 1125:24]
  wire  controls_config_bready; // @[BFS.scala 1125:24]
  (*dont_touch = "true" *)reg [31:0] level; // @[BFS.scala 1126:22]
  (*dont_touch = "true" *)reg [2:0] status; // @[BFS.scala 1136:23]
  wire  start = controls_io_data_0[0] & ~controls_io_data_0[1]; // @[BFS.scala 1137:38]
  (*dont_touch = "true" *)reg  FIN_0; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_1; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_2; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_3; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_4; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_5; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_6; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_7; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_8; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_9; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_10; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_11; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_12; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_13; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_14; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_15; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_16; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_17; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_18; // @[BFS.scala 1138:20]
  (*dont_touch = "true" *)reg  FIN_19; // @[BFS.scala 1138:20]
  wire [63:0] _new_tep_T = {controls_io_data_12,controls_io_data_13}; // @[Cat.scala 30:58]
  wire [63:0] new_tep = _new_tep_T + io_traveled_edges; // @[BFS.scala 1139:65]
  reg [63:0] counterValue; // @[BFS.scala 1140:29]
  wire  _controls_io_writeFlag_0_T = status == 3'h3; // @[BFS.scala 1143:38]
  wire  _controls_io_writeFlag_0_T_1 = status == 3'h2; // @[BFS.scala 1143:59]
  wire  _controls_io_writeFlag_0_T_3 = status == 3'h2 & io_signal_ack; // @[BFS.scala 1143:70]
  wire  _controls_io_writeFlag_0_T_5 = status == 3'h6; // @[BFS.scala 1143:108]
  wire [3:0] _controls_io_wptr_0_T_3 = _controls_io_writeFlag_0_T_1 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_0_T_4 = _controls_io_writeFlag_0_T_5 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_0_T_6 = _controls_io_wptr_0_T_3 | _controls_io_wptr_0_T_4; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_5 = _controls_io_writeFlag_0_T_1 ? new_tep[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_6 = _controls_io_writeFlag_0_T_5 ? counterValue[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [1:0] _controls_io_dataIn_0_T_7 = _controls_io_writeFlag_0_T ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_8 = _controls_io_dataIn_0_T_5 | _controls_io_dataIn_0_T_6; // @[Mux.scala 27:72]
  wire [31:0] _GEN_52 = {{30'd0}, _controls_io_dataIn_0_T_7}; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_1_T_1 = _controls_io_writeFlag_0_T_1 ? 4'hd : 4'hf; // @[BFS.scala 1155:29]
  wire [31:0] _controls_io_dataIn_1_T_4 = _controls_io_writeFlag_0_T_1 ? new_tep[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_1_T_5 = _controls_io_writeFlag_0_T_5 ? counterValue[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1 = status == 3'h0 & start; // @[BFS.scala 1161:28]
  wire  _T_2 = status == 3'h4; // @[BFS.scala 1163:21]
  wire [2:0] _GEN_0 = io_data_28 == level ? 3'h6 : 3'h1; // @[BFS.scala 1168:44 BFS.scala 1169:14 BFS.scala 1171:14]
  wire [2:0] _GEN_1 = _controls_io_writeFlag_0_T_5 ? 3'h5 : status; // @[BFS.scala 1175:40 BFS.scala 1176:12 BFS.scala 1136:23]
  wire [2:0] _GEN_2 = status == 3'h5 & io_flush_cache_end ? 3'h3 : _GEN_1; // @[BFS.scala 1173:62 BFS.scala 1174:12]
  wire [2:0] _GEN_3 = _controls_io_writeFlag_0_T_3 ? _GEN_0 : _GEN_2; // @[BFS.scala 1167:60]
  wire  _GEN_7 = io_fin_0 | FIN_0; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_9 = io_fin_1 | FIN_1; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_11 = io_fin_2 | FIN_2; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_13 = io_fin_3 | FIN_3; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_15 = io_fin_4 | FIN_4; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_17 = io_fin_5 | FIN_5; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_19 = io_fin_6 | FIN_6; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_21 = io_fin_7 | FIN_7; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_23 = io_fin_8 | FIN_8; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_25 = io_fin_9 | FIN_9; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_27 = io_fin_10 | FIN_10; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_29 = io_fin_11 | FIN_11; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_31 = io_fin_12 | FIN_12; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_33 = io_fin_13 | FIN_13; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_35 = io_fin_14 | FIN_14; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_37 = io_fin_15 | FIN_15; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_39 = io_fin_16 | FIN_16; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_41 = io_fin_17 | FIN_17; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_43 = io_fin_18 | FIN_18; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire  _GEN_45 = io_fin_19 | FIN_19; // @[BFS.scala 1185:28 BFS.scala 1186:11 BFS.scala 1138:20]
  wire [31:0] _level_T_1 = level + 32'h1; // @[BFS.scala 1192:20]
  wire  global_start = _controls_io_writeFlag_0_T_3 & level == 32'hffffffff; // @[BFS.scala 1197:68]
  wire [63:0] _counterValue_T_1 = counterValue + 64'h1; // @[BFS.scala 1201:34]
  reg [63:0] performanceValue_0; // @[BFS.scala 1204:33]
  LookupTable controls ( // @[BFS.scala 1125:24]
    .clock(controls_clock),
    .reset(controls_reset),
    .io_data_0(controls_io_data_0),
    .io_data_1(controls_io_data_1),
    .io_data_2(controls_io_data_2),
    .io_data_3(controls_io_data_3),
    .io_data_4(controls_io_data_4),
    .io_data_7(controls_io_data_7),
    .io_data_12(controls_io_data_12),
    .io_data_13(controls_io_data_13),
    .io_data_16(controls_io_data_16),
    .io_data_17(controls_io_data_17),
    .io_data_18(controls_io_data_18),
    .io_data_19(controls_io_data_19),
    .io_data_20(controls_io_data_20),
    .io_data_21(controls_io_data_21),
    .io_data_22(controls_io_data_22),
    .io_data_23(controls_io_data_23),
    .io_data_24(controls_io_data_24),
    .io_data_25(controls_io_data_25),
    .io_data_26(controls_io_data_26),
    .io_data_27(controls_io_data_27),
    .io_data_28(controls_io_data_28),
    .io_data_29(controls_io_data_29),
    .io_dataIn_0(controls_io_dataIn_0),
    .io_dataIn_1(controls_io_dataIn_1),
    .io_writeFlag_0(controls_io_writeFlag_0),
    .io_writeFlag_1(controls_io_writeFlag_1),
    .io_wptr_0(controls_io_wptr_0),
    .io_wptr_1(controls_io_wptr_1),
    .config_awaddr(controls_config_awaddr),
    .config_awvalid(controls_config_awvalid),
    .config_awready(controls_config_awready),
    .config_araddr(controls_config_araddr),
    .config_arvalid(controls_config_arvalid),
    .config_arready(controls_config_arready),
    .config_wdata(controls_config_wdata),
    .config_wvalid(controls_config_wvalid),
    .config_wready(controls_config_wready),
    .config_rdata(controls_config_rdata),
    .config_rvalid(controls_config_rvalid),
    .config_rready(controls_config_rready),
    .config_bvalid(controls_config_bvalid),
    .config_bready(controls_config_bready)
  );
  assign io_data_0 = controls_io_data_0; // @[BFS.scala 1217:11]
  assign io_data_1 = controls_io_data_1; // @[BFS.scala 1217:11]
  assign io_data_2 = controls_io_data_2; // @[BFS.scala 1217:11]
  assign io_data_3 = controls_io_data_3; // @[BFS.scala 1217:11]
  assign io_data_4 = controls_io_data_4; // @[BFS.scala 1217:11]
  assign io_data_7 = controls_io_data_7; // @[BFS.scala 1217:11]
  assign io_data_16 = controls_io_data_16; // @[BFS.scala 1217:11]
  assign io_data_17 = controls_io_data_17; // @[BFS.scala 1217:11]
  assign io_data_18 = controls_io_data_18; // @[BFS.scala 1217:11]
  assign io_data_19 = controls_io_data_19; // @[BFS.scala 1217:11]
  assign io_data_20 = controls_io_data_20; // @[BFS.scala 1217:11]
  assign io_data_21 = controls_io_data_21; // @[BFS.scala 1217:11]
  assign io_data_22 = controls_io_data_22; // @[BFS.scala 1217:11]
  assign io_data_23 = controls_io_data_23; // @[BFS.scala 1217:11]
  assign io_data_24 = controls_io_data_24; // @[BFS.scala 1217:11]
  assign io_data_25 = controls_io_data_25; // @[BFS.scala 1217:11]
  assign io_data_26 = controls_io_data_26; // @[BFS.scala 1217:11]
  assign io_data_27 = controls_io_data_27; // @[BFS.scala 1217:11]
  assign io_data_28 = controls_io_data_28; // @[BFS.scala 1217:11]
  assign io_data_29 = controls_io_data_29; // @[BFS.scala 1217:11]
  assign io_signal = _T_2 | _controls_io_writeFlag_0_T_1 & io_data_28 != level; // @[BFS.scala 1216:36]
  assign io_start = status == 3'h4; // @[BFS.scala 1219:22]
  assign io_level = level; // @[BFS.scala 1218:12]
  assign io_config_awready = controls_config_awready; // @[BFS.scala 1142:19]
  assign io_config_arready = controls_config_arready; // @[BFS.scala 1142:19]
  assign io_config_wready = controls_config_wready; // @[BFS.scala 1142:19]
  assign io_config_rdata = controls_config_rdata; // @[BFS.scala 1142:19]
  assign io_config_rvalid = controls_config_rvalid; // @[BFS.scala 1142:19]
  assign io_config_bvalid = controls_config_bvalid; // @[BFS.scala 1142:19]
  assign io_flush_cache = status == 3'h5; // @[BFS.scala 1220:28]
  assign controls_clock = clock;
  assign controls_reset = reset;
  assign controls_io_dataIn_0 = _controls_io_dataIn_0_T_8 | _GEN_52; // @[Mux.scala 27:72]
  assign controls_io_dataIn_1 = _controls_io_dataIn_1_T_4 | _controls_io_dataIn_1_T_5; // @[Mux.scala 27:72]
  assign controls_io_writeFlag_0 = status == 3'h3 | status == 3'h2 & io_signal_ack | status == 3'h6; // @[BFS.scala 1143:99]
  assign controls_io_writeFlag_1 = _controls_io_writeFlag_0_T_3 | _controls_io_writeFlag_0_T_5; // @[BFS.scala 1154:79]
  assign controls_io_wptr_0 = {{1'd0}, _controls_io_wptr_0_T_6}; // @[Mux.scala 27:72]
  assign controls_io_wptr_1 = {{1'd0}, _controls_io_wptr_1_T_1}; // @[BFS.scala 1155:29]
  assign controls_config_awaddr = io_config_awaddr; // @[BFS.scala 1142:19]
  assign controls_config_awvalid = io_config_awvalid; // @[BFS.scala 1142:19]
  assign controls_config_araddr = io_config_araddr; // @[BFS.scala 1142:19]
  assign controls_config_arvalid = io_config_arvalid; // @[BFS.scala 1142:19]
  assign controls_config_wdata = io_config_wdata; // @[BFS.scala 1142:19]
  assign controls_config_wvalid = io_config_wvalid; // @[BFS.scala 1142:19]
  assign controls_config_rready = io_config_rready; // @[BFS.scala 1142:19]
  assign controls_config_bready = io_config_bready; // @[BFS.scala 1142:19]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1126:22]
      level <= 32'h0; // @[BFS.scala 1126:22]
    end else if (_controls_io_writeFlag_0_T_3) begin // @[BFS.scala 1191:54]
      level <= _level_T_1; // @[BFS.scala 1192:11]
    end else if (_T_1) begin // @[BFS.scala 1193:43]
      level <= 32'hffffffff; // @[BFS.scala 1194:11]
    end
    if (reset) begin // @[BFS.scala 1136:23]
      status <= 3'h0; // @[BFS.scala 1136:23]
    end else if (status == 3'h0 & start) begin // @[BFS.scala 1161:37]
      status <= 3'h4; // @[BFS.scala 1162:12]
    end else if (status == 3'h4) begin // @[BFS.scala 1163:34]
      status <= 3'h1; // @[BFS.scala 1164:12]
    end else if (status == 3'h1 & (FIN_0 & FIN_1 & FIN_2 & FIN_3 & FIN_4 & FIN_5 & FIN_6 & FIN_7 & FIN_8 & FIN_9 &
      FIN_10 & FIN_11 & FIN_12 & FIN_13 & FIN_14 & FIN_15 & FIN_16 & FIN_17 & FIN_18 & FIN_19)) begin // @[BFS.scala 1165:51]
      status <= 3'h2; // @[BFS.scala 1166:12]
    end else begin
      status <= _GEN_3;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_0 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_0 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_0 <= _GEN_7;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_1 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_1 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_1 <= _GEN_9;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_2 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_2 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_2 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_3 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_3 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_3 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_4 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_4 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_4 <= _GEN_15;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_5 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_5 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_5 <= _GEN_17;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_6 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_6 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_6 <= _GEN_19;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_7 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_7 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_7 <= _GEN_21;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_8 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_8 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_8 <= _GEN_23;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_9 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_9 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_9 <= _GEN_25;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_10 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_10 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_10 <= _GEN_27;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_11 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_11 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_11 <= _GEN_29;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_12 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_12 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_12 <= _GEN_31;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_13 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_13 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_13 <= _GEN_33;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_14 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_14 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_14 <= _GEN_35;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_15 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_15 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_15 <= _GEN_37;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_16 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_16 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_16 <= _GEN_39;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_17 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_17 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_17 <= _GEN_41;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_18 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_18 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_18 <= _GEN_43;
    end
    if (reset) begin // @[BFS.scala 1138:20]
      FIN_19 <= 1'h0; // @[BFS.scala 1138:20]
    end else if (io_signal) begin // @[BFS.scala 1183:22]
      FIN_19 <= 1'h0; // @[BFS.scala 1184:11]
    end else begin
      FIN_19 <= _GEN_45;
    end
    if (reset) begin // @[BFS.scala 1140:29]
      counterValue <= 64'h0; // @[BFS.scala 1140:29]
    end else if (global_start) begin // @[BFS.scala 1198:22]
      counterValue <= 64'h0; // @[BFS.scala 1199:18]
    end else begin
      counterValue <= _counterValue_T_1; // @[BFS.scala 1201:18]
    end
    if (reset) begin // @[BFS.scala 1204:33]
      performanceValue_0 <= 64'h0; // @[BFS.scala 1204:33]
    end else if (global_start) begin // @[BFS.scala 1208:26]
      performanceValue_0 <= 64'h0; // @[BFS.scala 1209:29]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  level = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  status = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  FIN_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIN_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  FIN_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  FIN_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  FIN_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  FIN_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  FIN_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  FIN_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  FIN_8 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  FIN_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  FIN_10 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  FIN_11 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  FIN_12 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  FIN_13 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  FIN_14 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  FIN_15 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  FIN_16 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  FIN_17 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  FIN_18 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  FIN_19 = _RAND_21[0:0];
  _RAND_22 = {2{`RANDOM}};
  counterValue = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  performanceValue_0 = _RAND_23[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multi_port_mc(
  input          clock,
  input          reset,
  input          io_cacheable_out_ready,
  output         io_cacheable_out_valid,
  output [511:0] io_cacheable_out_bits_tdata,
  output [15:0]  io_cacheable_out_bits_tkeep,
  input  [31:0]  io_graph_scale,
  input          io_start,
  input          io_signal,
  input          io_end,
  output         io_signal_ack
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] tier_counter; // @[BFS.scala 1016:29]
  reg [31:0] tier_data_0; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_1; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_2; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_3; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_4; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_5; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_6; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_7; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_8; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_9; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_10; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_11; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_12; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_13; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_14; // @[BFS.scala 1017:26]
  reg [31:0] tier_data_15; // @[BFS.scala 1017:26]
  reg [2:0] status; // @[BFS.scala 1026:23]
  wire  _T = status == 3'h1; // @[BFS.scala 1030:19]
  wire  _T_2 = status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready; // @[BFS.scala 1030:67]
  wire [31:0] _tier_data_0_T_1 = tier_data_0 + 32'h40; // @[BFS.scala 1031:16]
  wire  _T_4 = io_signal & status == 3'h7; // @[BFS.scala 1032:28]
  wire [31:0] _tier_data_1_T_1 = tier_data_1 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_2_T_1 = tier_data_2 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_3_T_1 = tier_data_3 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_4_T_1 = tier_data_4 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_5_T_1 = tier_data_5 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_6_T_1 = tier_data_6 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_7_T_1 = tier_data_7 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_8_T_1 = tier_data_8 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_9_T_1 = tier_data_9 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_10_T_1 = tier_data_10 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_11_T_1 = tier_data_11 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_12_T_1 = tier_data_12 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_13_T_1 = tier_data_13 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_14_T_1 = tier_data_14 + 32'h40; // @[BFS.scala 1031:16]
  wire [31:0] _tier_data_15_T_1 = tier_data_15 + 32'h40; // @[BFS.scala 1031:16]
  wire  _T_81 = io_start & status == 3'h0; // @[BFS.scala 1038:17]
  wire [31:0] _tier_counter_T_2 = tier_counter - 32'h10; // @[BFS.scala 1041:59]
  wire  keep_0 = 32'h0 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_1 = 32'h1 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_2 = 32'h2 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_3 = 32'h3 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_4 = 32'h4 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_5 = 32'h5 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_6 = 32'h6 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_7 = 32'h7 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_8 = 32'h8 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_9 = 32'h9 < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_10 = 32'ha < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_11 = 32'hb < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_12 = 32'hc < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_13 = 32'hd < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_14 = 32'he < tier_counter; // @[BFS.scala 1045:52]
  wire  keep_15 = 32'hf < tier_counter; // @[BFS.scala 1045:52]
  wire  _T_94 = _T & tier_counter <= 32'h10 & tier_counter > 32'h0 & io_cacheable_out_valid; // @[BFS.scala 1049:89]
  wire  _T_96 = status == 3'h5; // @[BFS.scala 1052:21]
  wire [2:0] _GEN_35 = io_end ? 3'h0 : status; // @[BFS.scala 1056:21 BFS.scala 1057:12 BFS.scala 1026:23]
  wire [2:0] _GEN_36 = _T_4 ? 3'h1 : _GEN_35; // @[BFS.scala 1054:55 BFS.scala 1055:14]
  wire [255:0] io_cacheable_out_bits_tdata_lo = {tier_data_7,tier_data_6,tier_data_5,tier_data_4,tier_data_3,tier_data_2
    ,tier_data_1,tier_data_0}; // @[BFS.scala 1065:21]
  wire [511:0] _io_cacheable_out_bits_tdata_T_1 = {tier_data_15,tier_data_14,tier_data_13,tier_data_12,tier_data_11,
    tier_data_10,tier_data_9,tier_data_8,io_cacheable_out_bits_tdata_lo}; // @[BFS.scala 1065:21]
  wire [7:0] io_cacheable_out_bits_tkeep_lo = {keep_7,keep_6,keep_5,keep_4,keep_3,keep_2,keep_1,keep_0}; // @[BFS.scala 1066:87]
  wire [15:0] _io_cacheable_out_bits_tkeep_T_1 = {keep_15,keep_14,keep_13,keep_12,keep_11,keep_10,keep_9,keep_8,
    io_cacheable_out_bits_tkeep_lo}; // @[BFS.scala 1066:87]
  assign io_cacheable_out_valid = _T_96 | _T; // @[BFS.scala 1063:55]
  assign io_cacheable_out_bits_tdata = _T_96 ? 512'h80000000 : _io_cacheable_out_bits_tdata_T_1; // @[BFS.scala 1064:37]
  assign io_cacheable_out_bits_tkeep = _T_96 ? 16'h1 : _io_cacheable_out_bits_tkeep_T_1; // @[BFS.scala 1066:37]
  assign io_signal_ack = status == 3'h7; // @[BFS.scala 1083:27]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1016:29]
      tier_counter <= 32'h0; // @[BFS.scala 1016:29]
    end else if (io_start & status == 3'h0) begin // @[BFS.scala 1038:40]
      tier_counter <= io_graph_scale; // @[BFS.scala 1039:18]
    end else if (_T_2) begin // @[BFS.scala 1040:95]
      if (tier_counter > 32'h10) begin // @[BFS.scala 1041:24]
        tier_counter <= _tier_counter_T_2;
      end else begin
        tier_counter <= 32'h0;
      end
    end else if (_T_4) begin // @[BFS.scala 1042:55]
      tier_counter <= io_graph_scale; // @[BFS.scala 1043:18]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_0 <= 32'h0; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_0 <= _tier_data_0_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_0 <= 32'h0; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_1 <= 32'h4; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_1 <= _tier_data_1_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_1 <= 32'h4; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_2 <= 32'h8; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_2 <= _tier_data_2_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_2 <= 32'h8; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_3 <= 32'hc; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_3 <= _tier_data_3_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_3 <= 32'hc; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_4 <= 32'h10; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_4 <= _tier_data_4_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_4 <= 32'h10; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_5 <= 32'h14; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_5 <= _tier_data_5_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_5 <= 32'h14; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_6 <= 32'h18; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_6 <= _tier_data_6_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_6 <= 32'h18; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_7 <= 32'h1c; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_7 <= _tier_data_7_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_7 <= 32'h1c; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_8 <= 32'h20; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_8 <= _tier_data_8_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_8 <= 32'h20; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_9 <= 32'h24; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_9 <= _tier_data_9_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_9 <= 32'h24; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_10 <= 32'h28; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_10 <= _tier_data_10_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_10 <= 32'h28; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_11 <= 32'h2c; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_11 <= _tier_data_11_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_11 <= 32'h2c; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_12 <= 32'h30; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_12 <= _tier_data_12_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_12 <= 32'h30; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_13 <= 32'h34; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_13 <= _tier_data_13_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_13 <= 32'h34; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_14 <= 32'h38; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_14 <= _tier_data_14_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_14 <= 32'h38; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1017:26]
      tier_data_15 <= 32'h3c; // @[BFS.scala 1017:26]
    end else if (status == 3'h1 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1030:93]
      tier_data_15 <= _tier_data_15_T_1; // @[BFS.scala 1031:11]
    end else if (io_signal & status == 3'h7) begin // @[BFS.scala 1032:59]
      tier_data_15 <= 32'h3c; // @[BFS.scala 1033:11]
    end
    if (reset) begin // @[BFS.scala 1026:23]
      status <= 3'h0; // @[BFS.scala 1026:23]
    end else if (_T_81) begin // @[BFS.scala 1047:40]
      status <= 3'h1; // @[BFS.scala 1048:12]
    end else if (_T_94 & io_cacheable_out_ready) begin // @[BFS.scala 1050:54]
      status <= 3'h5; // @[BFS.scala 1051:12]
    end else if (status == 3'h5 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 1052:92]
      status <= 3'h7; // @[BFS.scala 1053:12]
    end else begin
      status <= _GEN_36;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tier_counter = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  tier_data_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  tier_data_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  tier_data_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  tier_data_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  tier_data_4 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  tier_data_5 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  tier_data_6 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  tier_data_7 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  tier_data_8 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  tier_data_9 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  tier_data_10 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  tier_data_11 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  tier_data_12 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  tier_data_13 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  tier_data_14 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  tier_data_15 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  status = _RAND_17[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_arbitrator(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  in_aclk; // @[util.scala 455:18]
  wire  in_aresetn; // @[util.scala 455:18]
  wire [511:0] in_s_axis_tdata; // @[util.scala 455:18]
  wire  in_s_axis_tvalid; // @[util.scala 455:18]
  wire [63:0] in_s_axis_tkeep; // @[util.scala 455:18]
  wire  in_s_axis_tready; // @[util.scala 455:18]
  wire  in_s_axis_tlast; // @[util.scala 455:18]
  wire [511:0] in_m_axis_tdata; // @[util.scala 455:18]
  wire  in_m_axis_tvalid; // @[util.scala 455:18]
  wire [63:0] in_m_axis_tkeep; // @[util.scala 455:18]
  wire  in_m_axis_tready; // @[util.scala 455:18]
  wire  in_m_axis_tlast; // @[util.scala 455:18]
  wire  mid_aclk; // @[util.scala 465:19]
  wire  mid_aresetn; // @[util.scala 465:19]
  wire [511:0] mid_s_axis_tdata; // @[util.scala 465:19]
  wire  mid_s_axis_tvalid; // @[util.scala 465:19]
  wire [63:0] mid_s_axis_tkeep; // @[util.scala 465:19]
  wire  mid_s_axis_tready; // @[util.scala 465:19]
  wire  mid_s_axis_tlast; // @[util.scala 465:19]
  wire [511:0] mid_m_axis_tdata; // @[util.scala 465:19]
  wire  mid_m_axis_tvalid; // @[util.scala 465:19]
  wire [63:0] mid_m_axis_tkeep; // @[util.scala 465:19]
  wire  mid_m_axis_tready; // @[util.scala 465:19]
  wire  mid_m_axis_tlast; // @[util.scala 465:19]
  wire  out_aclk; // @[util.scala 485:19]
  wire  out_aresetn; // @[util.scala 485:19]
  wire [31:0] out_s_axis_tdata; // @[util.scala 485:19]
  wire  out_s_axis_tvalid; // @[util.scala 485:19]
  wire [3:0] out_s_axis_tkeep; // @[util.scala 485:19]
  wire  out_s_axis_tready; // @[util.scala 485:19]
  wire  out_s_axis_tlast; // @[util.scala 485:19]
  wire [31:0] out_m_axis_tdata; // @[util.scala 485:19]
  wire  out_m_axis_tvalid; // @[util.scala 485:19]
  wire [3:0] out_m_axis_tkeep; // @[util.scala 485:19]
  wire  out_m_axis_tready; // @[util.scala 485:19]
  wire  out_m_axis_tlast; // @[util.scala 485:19]
  wire  in_keep_0 = in_m_axis_tkeep[0]; // @[util.scala 463:97]
  wire  in_keep_1 = in_m_axis_tkeep[1]; // @[util.scala 463:97]
  wire  in_keep_2 = in_m_axis_tkeep[2]; // @[util.scala 463:97]
  wire  in_keep_3 = in_m_axis_tkeep[3]; // @[util.scala 463:97]
  wire  in_keep_4 = in_m_axis_tkeep[4]; // @[util.scala 463:97]
  wire  in_keep_5 = in_m_axis_tkeep[5]; // @[util.scala 463:97]
  wire  in_keep_6 = in_m_axis_tkeep[6]; // @[util.scala 463:97]
  wire  in_keep_7 = in_m_axis_tkeep[7]; // @[util.scala 463:97]
  wire  in_keep_8 = in_m_axis_tkeep[8]; // @[util.scala 463:97]
  wire  in_keep_9 = in_m_axis_tkeep[9]; // @[util.scala 463:97]
  wire  in_keep_10 = in_m_axis_tkeep[10]; // @[util.scala 463:97]
  wire  in_keep_11 = in_m_axis_tkeep[11]; // @[util.scala 463:97]
  wire  in_keep_12 = in_m_axis_tkeep[12]; // @[util.scala 463:97]
  wire  in_keep_13 = in_m_axis_tkeep[13]; // @[util.scala 463:97]
  wire  in_keep_14 = in_m_axis_tkeep[14]; // @[util.scala 463:97]
  wire  in_keep_15 = in_m_axis_tkeep[15]; // @[util.scala 463:97]
  wire [4:0] _in_count_WIRE = {{4'd0}, in_keep_0}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_WIRE_1 = {{4'd0}, in_keep_1}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_1 = _in_count_WIRE + _in_count_WIRE_1; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_2 = {{4'd0}, in_keep_2}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_3 = _in_count_T_1 + _in_count_WIRE_2; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_3 = {{4'd0}, in_keep_3}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_5 = _in_count_T_3 + _in_count_WIRE_3; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_4 = {{4'd0}, in_keep_4}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_7 = _in_count_T_5 + _in_count_WIRE_4; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_5 = {{4'd0}, in_keep_5}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_9 = _in_count_T_7 + _in_count_WIRE_5; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_6 = {{4'd0}, in_keep_6}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_11 = _in_count_T_9 + _in_count_WIRE_6; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_7 = {{4'd0}, in_keep_7}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_13 = _in_count_T_11 + _in_count_WIRE_7; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_8 = {{4'd0}, in_keep_8}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_15 = _in_count_T_13 + _in_count_WIRE_8; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_9 = {{4'd0}, in_keep_9}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_17 = _in_count_T_15 + _in_count_WIRE_9; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_10 = {{4'd0}, in_keep_10}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_19 = _in_count_T_17 + _in_count_WIRE_10; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_11 = {{4'd0}, in_keep_11}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_21 = _in_count_T_19 + _in_count_WIRE_11; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_12 = {{4'd0}, in_keep_12}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_23 = _in_count_T_21 + _in_count_WIRE_12; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_13 = {{4'd0}, in_keep_13}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_25 = _in_count_T_23 + _in_count_WIRE_13; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_14 = {{4'd0}, in_keep_14}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] _in_count_T_27 = _in_count_T_25 + _in_count_WIRE_14; // @[util.scala 464:82]
  wire [4:0] _in_count_WIRE_15 = {{4'd0}, in_keep_15}; // @[util.scala 464:43 util.scala 464:43]
  wire [4:0] in_count = _in_count_T_27 + _in_count_WIRE_15; // @[util.scala 464:82]
  wire [58:0] mid_io_s_axis_tkeep_lo = in_m_axis_tkeep[58:0]; // @[util.scala 472:58]
  wire  keep_0 = mid_m_axis_tkeep[0]; // @[util.scala 476:95]
  wire  keep_1 = mid_m_axis_tkeep[1]; // @[util.scala 476:95]
  wire  keep_2 = mid_m_axis_tkeep[2]; // @[util.scala 476:95]
  wire  keep_3 = mid_m_axis_tkeep[3]; // @[util.scala 476:95]
  wire  keep_4 = mid_m_axis_tkeep[4]; // @[util.scala 476:95]
  wire  keep_5 = mid_m_axis_tkeep[5]; // @[util.scala 476:95]
  wire  keep_6 = mid_m_axis_tkeep[6]; // @[util.scala 476:95]
  wire  keep_7 = mid_m_axis_tkeep[7]; // @[util.scala 476:95]
  wire  keep_8 = mid_m_axis_tkeep[8]; // @[util.scala 476:95]
  wire  keep_9 = mid_m_axis_tkeep[9]; // @[util.scala 476:95]
  wire  keep_10 = mid_m_axis_tkeep[10]; // @[util.scala 476:95]
  wire  keep_11 = mid_m_axis_tkeep[11]; // @[util.scala 476:95]
  wire  keep_12 = mid_m_axis_tkeep[12]; // @[util.scala 476:95]
  wire  keep_13 = mid_m_axis_tkeep[13]; // @[util.scala 476:95]
  wire  keep_14 = mid_m_axis_tkeep[14]; // @[util.scala 476:95]
  wire  keep_15 = mid_m_axis_tkeep[15]; // @[util.scala 476:95]
  reg  index_0; // @[util.scala 477:22]
  reg  index_1; // @[util.scala 477:22]
  reg  index_2; // @[util.scala 477:22]
  reg  index_3; // @[util.scala 477:22]
  reg  index_4; // @[util.scala 477:22]
  reg  index_5; // @[util.scala 477:22]
  reg  index_6; // @[util.scala 477:22]
  reg  index_7; // @[util.scala 477:22]
  reg  index_8; // @[util.scala 477:22]
  reg  index_9; // @[util.scala 477:22]
  reg  index_10; // @[util.scala 477:22]
  reg  index_11; // @[util.scala 477:22]
  reg  index_12; // @[util.scala 477:22]
  reg  index_13; // @[util.scala 477:22]
  reg  index_14; // @[util.scala 477:22]
  reg  index_15; // @[util.scala 477:22]
  wire  ungrant_keep_0 = keep_0 & ~index_0; // @[util.scala 479:22]
  wire  ungrant_keep_1 = keep_1 & ~index_1; // @[util.scala 479:22]
  wire  ungrant_keep_2 = keep_2 & ~index_2; // @[util.scala 479:22]
  wire  ungrant_keep_3 = keep_3 & ~index_3; // @[util.scala 479:22]
  wire  ungrant_keep_4 = keep_4 & ~index_4; // @[util.scala 479:22]
  wire  ungrant_keep_5 = keep_5 & ~index_5; // @[util.scala 479:22]
  wire  ungrant_keep_6 = keep_6 & ~index_6; // @[util.scala 479:22]
  wire  ungrant_keep_7 = keep_7 & ~index_7; // @[util.scala 479:22]
  wire  ungrant_keep_8 = keep_8 & ~index_8; // @[util.scala 479:22]
  wire  ungrant_keep_9 = keep_9 & ~index_9; // @[util.scala 479:22]
  wire  ungrant_keep_10 = keep_10 & ~index_10; // @[util.scala 479:22]
  wire  ungrant_keep_11 = keep_11 & ~index_11; // @[util.scala 479:22]
  wire  ungrant_keep_12 = keep_12 & ~index_12; // @[util.scala 479:22]
  wire  ungrant_keep_13 = keep_13 & ~index_13; // @[util.scala 479:22]
  wire  ungrant_keep_14 = keep_14 & ~index_14; // @[util.scala 479:22]
  wire  ungrant_keep_15 = keep_15 & ~index_15; // @[util.scala 479:22]
  wire  grant_1 = ~ungrant_keep_0; // @[util.scala 363:78]
  wire  grant_2 = ~(ungrant_keep_0 | ungrant_keep_1); // @[util.scala 363:78]
  wire  grant_3 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2); // @[util.scala 363:78]
  wire  grant_4 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3); // @[util.scala 363:78]
  wire  grant_5 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4); // @[util.scala 363:78]
  wire  grant_6 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5)
    ; // @[util.scala 363:78]
  wire  grant_7 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6); // @[util.scala 363:78]
  wire  grant_8 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7); // @[util.scala 363:78]
  wire  grant_9 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8); // @[util.scala 363:78]
  wire  grant_10 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9); // @[util.scala 363:78]
  wire  grant_11 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10); // @[util.scala 363:78]
  wire  grant_12 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10 | ungrant_keep_11); // @[util.scala 363:78]
  wire  grant_13 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10 | ungrant_keep_11 |
    ungrant_keep_12); // @[util.scala 363:78]
  wire  grant_14 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10 | ungrant_keep_11 |
    ungrant_keep_12 | ungrant_keep_13); // @[util.scala 363:78]
  wire  grant_15 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2 | ungrant_keep_3 | ungrant_keep_4 | ungrant_keep_5
     | ungrant_keep_6 | ungrant_keep_7 | ungrant_keep_8 | ungrant_keep_9 | ungrant_keep_10 | ungrant_keep_11 |
    ungrant_keep_12 | ungrant_keep_13 | ungrant_keep_14); // @[util.scala 363:78]
  wire  choosen_keep_1 = grant_1 & ungrant_keep_1; // @[util.scala 483:22]
  wire  choosen_keep_2 = grant_2 & ungrant_keep_2; // @[util.scala 483:22]
  wire  choosen_keep_3 = grant_3 & ungrant_keep_3; // @[util.scala 483:22]
  wire  choosen_keep_4 = grant_4 & ungrant_keep_4; // @[util.scala 483:22]
  wire  choosen_keep_5 = grant_5 & ungrant_keep_5; // @[util.scala 483:22]
  wire  choosen_keep_6 = grant_6 & ungrant_keep_6; // @[util.scala 483:22]
  wire  choosen_keep_7 = grant_7 & ungrant_keep_7; // @[util.scala 483:22]
  wire  choosen_keep_8 = grant_8 & ungrant_keep_8; // @[util.scala 483:22]
  wire  choosen_keep_9 = grant_9 & ungrant_keep_9; // @[util.scala 483:22]
  wire  choosen_keep_10 = grant_10 & ungrant_keep_10; // @[util.scala 483:22]
  wire  choosen_keep_11 = grant_11 & ungrant_keep_11; // @[util.scala 483:22]
  wire  choosen_keep_12 = grant_12 & ungrant_keep_12; // @[util.scala 483:22]
  wire  choosen_keep_13 = grant_13 & ungrant_keep_13; // @[util.scala 483:22]
  wire  choosen_keep_14 = grant_14 & ungrant_keep_14; // @[util.scala 483:22]
  wire  choosen_keep_15 = grant_15 & ungrant_keep_15; // @[util.scala 483:22]
  wire  _T_1 = mid_m_axis_tvalid; // @[util.scala 491:72]
  wire  _T_4 = out_s_axis_tready; // @[util.scala 493:78]
  wire  _T_5 = out_s_axis_tvalid & out_s_axis_tready; // @[util.scala 493:48]
  reg [4:0] count; // @[util.scala 499:22]
  wire [4:0] next_count = mid_m_axis_tkeep[63:59]; // @[util.scala 500:39]
  wire [4:0] _count_T_1 = next_count - 5'h1; // @[util.scala 503:27]
  wire [4:0] _count_T_3 = count - 5'h1; // @[util.scala 505:22]
  wire [31:0] _out_io_s_axis_tdata_T_16 = ungrant_keep_0 ? mid_m_axis_tdata[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_17 = choosen_keep_1 ? mid_m_axis_tdata[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_18 = choosen_keep_2 ? mid_m_axis_tdata[95:64] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_19 = choosen_keep_3 ? mid_m_axis_tdata[127:96] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_20 = choosen_keep_4 ? mid_m_axis_tdata[159:128] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_21 = choosen_keep_5 ? mid_m_axis_tdata[191:160] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_22 = choosen_keep_6 ? mid_m_axis_tdata[223:192] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_23 = choosen_keep_7 ? mid_m_axis_tdata[255:224] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_24 = choosen_keep_8 ? mid_m_axis_tdata[287:256] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_25 = choosen_keep_9 ? mid_m_axis_tdata[319:288] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_26 = choosen_keep_10 ? mid_m_axis_tdata[351:320] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_27 = choosen_keep_11 ? mid_m_axis_tdata[383:352] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_28 = choosen_keep_12 ? mid_m_axis_tdata[415:384] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_29 = choosen_keep_13 ? mid_m_axis_tdata[447:416] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_30 = choosen_keep_14 ? mid_m_axis_tdata[479:448] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_31 = choosen_keep_15 ? mid_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_32 = _out_io_s_axis_tdata_T_16 | _out_io_s_axis_tdata_T_17; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_33 = _out_io_s_axis_tdata_T_32 | _out_io_s_axis_tdata_T_18; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_34 = _out_io_s_axis_tdata_T_33 | _out_io_s_axis_tdata_T_19; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_35 = _out_io_s_axis_tdata_T_34 | _out_io_s_axis_tdata_T_20; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_36 = _out_io_s_axis_tdata_T_35 | _out_io_s_axis_tdata_T_21; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_37 = _out_io_s_axis_tdata_T_36 | _out_io_s_axis_tdata_T_22; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_38 = _out_io_s_axis_tdata_T_37 | _out_io_s_axis_tdata_T_23; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_39 = _out_io_s_axis_tdata_T_38 | _out_io_s_axis_tdata_T_24; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_40 = _out_io_s_axis_tdata_T_39 | _out_io_s_axis_tdata_T_25; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_41 = _out_io_s_axis_tdata_T_40 | _out_io_s_axis_tdata_T_26; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_42 = _out_io_s_axis_tdata_T_41 | _out_io_s_axis_tdata_T_27; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_43 = _out_io_s_axis_tdata_T_42 | _out_io_s_axis_tdata_T_28; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_44 = _out_io_s_axis_tdata_T_43 | _out_io_s_axis_tdata_T_29; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_45 = _out_io_s_axis_tdata_T_44 | _out_io_s_axis_tdata_T_30; // @[Mux.scala 27:72]
  axis_arbitrator_in_reg_slice_64 in ( // @[util.scala 455:18]
    .aclk(in_aclk),
    .aresetn(in_aresetn),
    .s_axis_tdata(in_s_axis_tdata),
    .s_axis_tvalid(in_s_axis_tvalid),
    .s_axis_tkeep(in_s_axis_tkeep),
    .s_axis_tready(in_s_axis_tready),
    .s_axis_tlast(in_s_axis_tlast),
    .m_axis_tdata(in_m_axis_tdata),
    .m_axis_tvalid(in_m_axis_tvalid),
    .m_axis_tkeep(in_m_axis_tkeep),
    .m_axis_tready(in_m_axis_tready),
    .m_axis_tlast(in_m_axis_tlast)
  );
  axis_arbitrator_in_reg_slice_64 mid ( // @[util.scala 465:19]
    .aclk(mid_aclk),
    .aresetn(mid_aresetn),
    .s_axis_tdata(mid_s_axis_tdata),
    .s_axis_tvalid(mid_s_axis_tvalid),
    .s_axis_tkeep(mid_s_axis_tkeep),
    .s_axis_tready(mid_s_axis_tready),
    .s_axis_tlast(mid_s_axis_tlast),
    .m_axis_tdata(mid_m_axis_tdata),
    .m_axis_tvalid(mid_m_axis_tvalid),
    .m_axis_tkeep(mid_m_axis_tkeep),
    .m_axis_tready(mid_m_axis_tready),
    .m_axis_tlast(mid_m_axis_tlast)
  );
  axis_arbitrator_out_reg_slice_4 out ( // @[util.scala 485:19]
    .aclk(out_aclk),
    .aresetn(out_aresetn),
    .s_axis_tdata(out_s_axis_tdata),
    .s_axis_tvalid(out_s_axis_tvalid),
    .s_axis_tkeep(out_s_axis_tkeep),
    .s_axis_tready(out_s_axis_tready),
    .s_axis_tlast(out_s_axis_tlast),
    .m_axis_tdata(out_m_axis_tdata),
    .m_axis_tvalid(out_m_axis_tvalid),
    .m_axis_tkeep(out_m_axis_tkeep),
    .m_axis_tready(out_m_axis_tready),
    .m_axis_tlast(out_m_axis_tlast)
  );
  assign io_xbar_in_ready = in_s_axis_tready; // @[util.scala 461:20]
  assign io_ddr_out_valid = out_m_axis_tvalid; // @[util.scala 516:20]
  assign io_ddr_out_bits_tdata = out_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign in_aclk = clock; // @[util.scala 457:29]
  assign in_aresetn = ~reset; // @[util.scala 458:20]
  assign in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_s_axis_tvalid = io_xbar_in_valid; // @[util.scala 460:23]
  assign in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign in_m_axis_tready = mid_s_axis_tready; // @[util.scala 473:23]
  assign mid_aclk = clock; // @[util.scala 467:30]
  assign mid_aresetn = ~reset; // @[util.scala 468:21]
  assign mid_s_axis_tdata = in_m_axis_tdata; // @[util.scala 470:23]
  assign mid_s_axis_tvalid = in_m_axis_tvalid; // @[util.scala 469:24]
  assign mid_s_axis_tkeep = {in_count,mid_io_s_axis_tkeep_lo}; // @[Cat.scala 30:58]
  assign mid_s_axis_tlast = in_m_axis_tlast; // @[util.scala 471:23]
  assign mid_m_axis_tready = _T_4 & (count == 5'h1 | next_count == 5'h1); // @[util.scala 508:57]
  assign out_aclk = clock; // @[util.scala 486:30]
  assign out_aresetn = ~reset; // @[util.scala 487:21]
  assign out_s_axis_tdata = _out_io_s_axis_tdata_T_45 | _out_io_s_axis_tdata_T_31; // @[Mux.scala 27:72]
  assign out_s_axis_tvalid = (ungrant_keep_0 | choosen_keep_1 | choosen_keep_2 | choosen_keep_3 | choosen_keep_4 |
    choosen_keep_5 | choosen_keep_6 | choosen_keep_7 | choosen_keep_8 | choosen_keep_9 | choosen_keep_10 |
    choosen_keep_11 | choosen_keep_12 | choosen_keep_13 | choosen_keep_14 | choosen_keep_15) & _T_1; // @[util.scala 510:52]
  assign out_s_axis_tkeep = 4'h1; // @[util.scala 511:23]
  assign out_s_axis_tlast = 1'h1; // @[util.scala 512:23]
  assign out_m_axis_tready = io_ddr_out_ready; // @[util.scala 517:24]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 477:22]
      index_0 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_0 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_0 <= index_0 | ungrant_keep_0; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_1 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_1 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_1 <= index_1 | choosen_keep_1; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_2 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_2 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_2 <= index_2 | choosen_keep_2; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_3 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_3 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_3 <= index_3 | choosen_keep_3; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_4 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_4 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_4 <= index_4 | choosen_keep_4; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_5 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_5 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_5 <= index_5 | choosen_keep_5; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_6 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_6 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_6 <= index_6 | choosen_keep_6; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_7 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_7 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_7 <= index_7 | choosen_keep_7; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_8 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_8 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_8 <= index_8 | choosen_keep_8; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_9 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_9 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_9 <= index_9 | choosen_keep_9; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_10 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_10 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_10 <= index_10 | choosen_keep_10; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_11 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_11 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_11 <= index_11 | choosen_keep_11; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_12 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_12 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_12 <= index_12 | choosen_keep_12; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_13 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_13 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_13 <= index_13 | choosen_keep_13; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_14 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_14 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_14 <= index_14 | choosen_keep_14; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_15 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_15 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_15 <= index_15 | choosen_keep_15; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 499:22]
      count <= 5'h0; // @[util.scala 499:22]
    end else if (_T_5) begin // @[util.scala 501:71]
      if (count == 5'h0) begin // @[util.scala 502:24]
        count <= _count_T_1; // @[util.scala 503:13]
      end else begin
        count <= _count_T_3; // @[util.scala 505:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  index_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  index_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  index_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  index_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  index_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  index_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  index_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  index_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  index_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  index_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  index_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  index_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  index_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  index_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  index_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  index_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  count = _RAND_16[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h0 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h0 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h0 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h0 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h0 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h0 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h0 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h0 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h0 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h0 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h0 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h0 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h0 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h0 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h0 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h0 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  (*dont_touch = "true" *)reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  (*dont_touch = "true" *)reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_1(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h1 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h1 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h1 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h1 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h1 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h1 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h1 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h1 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h1 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h1 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h1 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h1 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h1 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h1 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h1 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h1 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_2(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h2 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h2 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h2 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h2 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h2 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h2 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h2 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h2 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h2 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h2 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h2 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h2 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h2 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h2 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h2 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h2 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_3(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h3 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h3 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h3 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h3 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h3 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h3 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h3 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h3 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h3 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h3 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h3 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h3 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h3 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h3 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h3 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h3 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_4(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h4 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h4 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h4 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h4 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h4 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h4 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h4 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h4 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h4 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h4 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h4 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h4 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h4 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h4 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h4 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h4 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_5(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h5 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h5 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h5 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h5 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h5 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h5 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h5 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h5 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h5 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h5 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h5 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h5 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h5 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h5 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h5 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h5 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_6(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h6 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h6 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h6 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h6 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h6 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h6 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h6 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h6 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h6 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h6 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h6 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h6 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h6 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h6 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h6 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h6 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_7(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h7 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h7 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h7 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h7 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h7 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h7 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h7 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h7 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h7 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h7 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h7 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h7 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h7 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h7 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h7 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h7 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_8(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h8 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h8 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h8 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h8 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h8 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h8 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h8 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h8 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h8 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h8 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h8 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h8 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h8 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h8 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h8 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h8 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_9(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'h9 & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'h9 & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'h9 & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'h9 & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'h9 & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'h9 & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'h9 & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'h9 & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'h9 & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'h9 & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'h9 & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'h9 & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'h9 & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'h9 & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'h9 & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'h9 & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_10(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'ha & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'ha & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'ha & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'ha & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'ha & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'ha & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'ha & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'ha & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'ha & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'ha & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'ha & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'ha & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'ha & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'ha & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'ha & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'ha & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_11(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'hb & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'hb & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'hb & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'hb & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'hb & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'hb & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'hb & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'hb & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'hb & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'hb & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'hb & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'hb & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'hb & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'hb & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'hb & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'hb & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_12(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'hc & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'hc & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'hc & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'hc & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'hc & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'hc & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'hc & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'hc & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'hc & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'hc & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'hc & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'hc & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'hc & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'hc & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'hc & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'hc & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_13(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'hd & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'hd & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'hd & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'hd & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'hd & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'hd & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'hd & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'hd & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'hd & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'hd & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'hd & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'hd & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'hd & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'hd & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'hd & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'hd & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_14(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'he & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'he & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'he & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'he & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'he & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'he & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'he & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'he & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'he & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'he & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'he & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'he & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'he & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'he & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'he & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'he & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter_15(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  output         io_end,
  input  [2:0]   io_local_fpga_id,
  input  [31:0]  io_graph_scale
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] bitmap__addra; // @[BFS.scala 802:22]
  wire  bitmap__clka; // @[BFS.scala 802:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 802:22]
  wire  bitmap__ena; // @[BFS.scala 802:22]
  wire  bitmap__wea; // @[BFS.scala 802:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 802:22]
  wire  bitmap__clkb; // @[BFS.scala 802:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 802:22]
  wire  bitmap__enb; // @[BFS.scala 802:22]
  wire  arbi_clock; // @[BFS.scala 803:20]
  wire  arbi_reset; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 803:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 803:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 803:20]
  wire  arbi_io_xbar_in_bits_tlast; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 803:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 803:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 803:20]
  wire  scatter_in_aclk; // @[BFS.scala 828:26]
  wire  scatter_in_aresetn; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_s_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_s_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_s_axis_tlast; // @[BFS.scala 828:26]
  wire [511:0] scatter_in_m_axis_tdata; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tvalid; // @[BFS.scala 828:26]
  wire [63:0] scatter_in_m_axis_tkeep; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tready; // @[BFS.scala 828:26]
  wire  scatter_in_m_axis_tlast; // @[BFS.scala 828:26]
  wire  vertex_in_fifo_s_axis_aclk; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_s_axis_tid; // @[BFS.scala 844:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 844:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tready; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[BFS.scala 844:30]
  wire  vertex_in_fifo_m_axis_tid; // @[BFS.scala 844:30]
  wire  vertex_out_fifo_aclk; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_aresetn; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 857:31]
  wire [31:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 857:31]
  wire [3:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 857:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 857:31]
  reg [2:0] local_fpga_id; // @[BFS.scala 804:30]
  wire [2:0] _GEN_13 = {{1'd0}, scatter_in_m_axis_tdata[1:0]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_6 = _GEN_13 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_0_T_7 = scatter_in_m_axis_tdata[5:2] == 4'hf & _filtered_keep_0_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_0_T_8 = scatter_in_m_axis_tdata[31] | _filtered_keep_0_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_0 = scatter_in_m_axis_tkeep[0] & _filtered_keep_0_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_14 = {{1'd0}, scatter_in_m_axis_tdata[33:32]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_6 = _GEN_14 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_1_T_7 = scatter_in_m_axis_tdata[37:34] == 4'hf & _filtered_keep_1_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_1_T_8 = scatter_in_m_axis_tdata[63] | _filtered_keep_1_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_1 = scatter_in_m_axis_tkeep[1] & _filtered_keep_1_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_15 = {{1'd0}, scatter_in_m_axis_tdata[65:64]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_6 = _GEN_15 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_2_T_7 = scatter_in_m_axis_tdata[69:66] == 4'hf & _filtered_keep_2_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_2_T_8 = scatter_in_m_axis_tdata[95] | _filtered_keep_2_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_2 = scatter_in_m_axis_tkeep[2] & _filtered_keep_2_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_16 = {{1'd0}, scatter_in_m_axis_tdata[97:96]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_6 = _GEN_16 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_3_T_7 = scatter_in_m_axis_tdata[101:98] == 4'hf & _filtered_keep_3_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_3_T_8 = scatter_in_m_axis_tdata[127] | _filtered_keep_3_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_3 = scatter_in_m_axis_tkeep[3] & _filtered_keep_3_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_17 = {{1'd0}, scatter_in_m_axis_tdata[129:128]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_6 = _GEN_17 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_4_T_7 = scatter_in_m_axis_tdata[133:130] == 4'hf & _filtered_keep_4_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_4_T_8 = scatter_in_m_axis_tdata[159] | _filtered_keep_4_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_4 = scatter_in_m_axis_tkeep[4] & _filtered_keep_4_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_18 = {{1'd0}, scatter_in_m_axis_tdata[161:160]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_6 = _GEN_18 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_5_T_7 = scatter_in_m_axis_tdata[165:162] == 4'hf & _filtered_keep_5_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_5_T_8 = scatter_in_m_axis_tdata[191] | _filtered_keep_5_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_5 = scatter_in_m_axis_tkeep[5] & _filtered_keep_5_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_19 = {{1'd0}, scatter_in_m_axis_tdata[193:192]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_6 = _GEN_19 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_6_T_7 = scatter_in_m_axis_tdata[197:194] == 4'hf & _filtered_keep_6_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_6_T_8 = scatter_in_m_axis_tdata[223] | _filtered_keep_6_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_6 = scatter_in_m_axis_tkeep[6] & _filtered_keep_6_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_20 = {{1'd0}, scatter_in_m_axis_tdata[225:224]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_6 = _GEN_20 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_7_T_7 = scatter_in_m_axis_tdata[229:226] == 4'hf & _filtered_keep_7_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_7_T_8 = scatter_in_m_axis_tdata[255] | _filtered_keep_7_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_7 = scatter_in_m_axis_tkeep[7] & _filtered_keep_7_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_21 = {{1'd0}, scatter_in_m_axis_tdata[257:256]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_6 = _GEN_21 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_8_T_7 = scatter_in_m_axis_tdata[261:258] == 4'hf & _filtered_keep_8_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_8_T_8 = scatter_in_m_axis_tdata[287] | _filtered_keep_8_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_8 = scatter_in_m_axis_tkeep[8] & _filtered_keep_8_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_22 = {{1'd0}, scatter_in_m_axis_tdata[289:288]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_6 = _GEN_22 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_9_T_7 = scatter_in_m_axis_tdata[293:290] == 4'hf & _filtered_keep_9_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_9_T_8 = scatter_in_m_axis_tdata[319] | _filtered_keep_9_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_9 = scatter_in_m_axis_tkeep[9] & _filtered_keep_9_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_23 = {{1'd0}, scatter_in_m_axis_tdata[321:320]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_6 = _GEN_23 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_10_T_7 = scatter_in_m_axis_tdata[325:322] == 4'hf & _filtered_keep_10_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_10_T_8 = scatter_in_m_axis_tdata[351] | _filtered_keep_10_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_10 = scatter_in_m_axis_tkeep[10] & _filtered_keep_10_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_24 = {{1'd0}, scatter_in_m_axis_tdata[353:352]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_6 = _GEN_24 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_11_T_7 = scatter_in_m_axis_tdata[357:354] == 4'hf & _filtered_keep_11_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_11_T_8 = scatter_in_m_axis_tdata[383] | _filtered_keep_11_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_11 = scatter_in_m_axis_tkeep[11] & _filtered_keep_11_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_25 = {{1'd0}, scatter_in_m_axis_tdata[385:384]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_6 = _GEN_25 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_12_T_7 = scatter_in_m_axis_tdata[389:386] == 4'hf & _filtered_keep_12_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_12_T_8 = scatter_in_m_axis_tdata[415] | _filtered_keep_12_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_12 = scatter_in_m_axis_tkeep[12] & _filtered_keep_12_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_26 = {{1'd0}, scatter_in_m_axis_tdata[417:416]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_6 = _GEN_26 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_13_T_7 = scatter_in_m_axis_tdata[421:418] == 4'hf & _filtered_keep_13_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_13_T_8 = scatter_in_m_axis_tdata[447] | _filtered_keep_13_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_13 = scatter_in_m_axis_tkeep[13] & _filtered_keep_13_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_27 = {{1'd0}, scatter_in_m_axis_tdata[449:448]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_6 = _GEN_27 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_14_T_7 = scatter_in_m_axis_tdata[453:450] == 4'hf & _filtered_keep_14_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_14_T_8 = scatter_in_m_axis_tdata[479] | _filtered_keep_14_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_14 = scatter_in_m_axis_tkeep[14] & _filtered_keep_14_T_8; // @[BFS.scala 838:15]
  wire [2:0] _GEN_28 = {{1'd0}, scatter_in_m_axis_tdata[481:480]}; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_6 = _GEN_28 == local_fpga_id; // @[BFS.scala 812:40]
  wire  _filtered_keep_15_T_7 = scatter_in_m_axis_tdata[485:482] == 4'hf & _filtered_keep_15_T_6; // @[BFS.scala 811:85]
  wire  _filtered_keep_15_T_8 = scatter_in_m_axis_tdata[511] | _filtered_keep_15_T_7; // @[BFS.scala 839:12]
  wire  filtered_keep_15 = scatter_in_m_axis_tkeep[15] & _filtered_keep_15_T_8; // @[BFS.scala 838:15]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 850:57]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[BFS.scala 850:57]
  wire [63:0] _arbi_io_xbar_in_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  halt = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 863:47]
  reg  bitmap_wait_valid; // @[BFS.scala 864:28]
  reg [31:0] bitmap_wait_bits; // @[BFS.scala 864:28]
  wire  _T = ~halt; // @[BFS.scala 865:8]
  reg  bitmap_write_addr_valid; // @[BFS.scala 870:34]
  reg [31:0] bitmap_write_addr_bits; // @[BFS.scala 870:34]
  wire [26:0] _GEN_29 = {{2'd0}, bitmap_wait_bits[30:6]}; // @[BFS.scala 823:59]
  wire  _bitmap_write_addr_valid_T_1 = _GEN_29 > 27'he7fff; // @[BFS.scala 823:59]
  wire [3:0] _bitmap_write_addr_valid_WIRE = {{1'd0}, bitmap_wait_bits[8:6]}; // @[BFS.scala 825:107 BFS.scala 825:107]
  wire [3:0] _bitmap_write_addr_valid_T_3 = _GEN_29 > 27'he7fff ? 4'h8 : _bitmap_write_addr_valid_WIRE; // @[BFS.scala 823:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_29 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE = {{5'd0}, bitmap_wait_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 817:8]
  wire [26:0] _GEN_32 = {{2'd0}, bitmap_write_addr_bits[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_32 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{5'd0}, bitmap_write_addr_bits[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_32 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 817:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 888:41]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_valid & bitmap_wait_valid & _bitmap_doutb_T_15; // @[BFS.scala 887:51]
  reg [8:0] bitmap_write_data_bits; // @[BFS.scala 876:34]
  reg  bitmap_write_data_forward_valid; // @[BFS.scala 882:42]
  reg [8:0] bitmap_write_data_forward_bits; // @[BFS.scala 882:42]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_valid ? bitmap_write_data_forward_bits : bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_valid_T_3; // @[BFS.scala 873:20]
  wire  _bitmap_write_addr_valid_T_9 = ~_bitmap_write_addr_valid_T_4[0] | bitmap_wait_bits[31]; // @[BFS.scala 873:71]
  wire [23:0] _bitmap_write_data_bits_T_4 = 24'h1 << _bitmap_write_addr_valid_T_3; // @[BFS.scala 880:56]
  wire [23:0] _GEN_36 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 880:44]
  wire [23:0] _bitmap_write_data_bits_T_5 = _GEN_36 | _bitmap_write_data_bits_T_4; // @[BFS.scala 880:44]
  wire [23:0] _GEN_5 = _T ? _bitmap_write_data_bits_T_5 : {{15'd0}, bitmap_write_data_bits}; // @[BFS.scala 877:14 BFS.scala 880:28 BFS.scala 876:34]
  wire [26:0] _GEN_37 = {{2'd0}, arbi_io_ddr_out_bits_tdata[30:6]}; // @[BFS.scala 817:59]
  wire [26:0] _bitmap_write_data_forward_valid_T_5 = _GEN_37 - 27'he7fff; // @[BFS.scala 818:57]
  wire [26:0] _bitmap_write_data_forward_valid_WIRE = {{5'd0}, arbi_io_ddr_out_bits_tdata[30:9]}; // @[BFS.scala 819:69 BFS.scala 819:69]
  wire [26:0] _bitmap_write_data_forward_valid_T_7 = _GEN_37 > 27'he7fff ? _bitmap_write_data_forward_valid_T_5 :
    _bitmap_write_data_forward_valid_WIRE; // @[BFS.scala 817:8]
  wire  _bitmap_write_data_forward_valid_T_15 = _bitmap_write_data_forward_valid_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 884:50]
  wire [26:0] _bitmap_io_addrb_T_14 = halt ? _bitmap_doutb_T_7 : _bitmap_write_data_forward_valid_T_7; // @[BFS.scala 894:25]
  reg [31:0] wb_bram; // @[BFS.scala 910:24]
  wire [31:0] aligned_graph_scale = {{19'd0}, io_graph_scale[31:19]}; // @[BFS.scala 912:45]
  reg [31:0] num_small_sp; // @[BFS.scala 914:29]
  wire [50:0] _GEN_48 = {aligned_graph_scale, 19'h0}; // @[BFS.scala 917:46]
  wire [62:0] _num_small_sp_T = {{12'd0}, _GEN_48}; // @[BFS.scala 917:46]
  wire [62:0] _GEN_49 = {{31'd0}, io_graph_scale}; // @[BFS.scala 917:23]
  wire  _num_small_sp_T_1 = _GEN_49 > _num_small_sp_T; // @[BFS.scala 917:23]
  wire [31:0] _GEN_50 = {{31'd0}, _num_small_sp_T_1}; // @[BFS.scala 916:41]
  wire [31:0] _num_small_sp_T_3 = aligned_graph_scale + _GEN_50; // @[BFS.scala 916:41]
  wire  _T_7 = wb_bram > 32'h0; // @[BFS.scala 918:22]
  wire  _T_9 = wb_bram > 32'h0 & wb_bram <= 32'h40; // @[BFS.scala 918:28]
  wire  _T_10 = num_small_sp != 32'h0; // @[BFS.scala 918:63]
  wire [31:0] _num_small_sp_T_5 = num_small_sp - 32'h1; // @[BFS.scala 919:34]
  wire  _vertices_per_sp_T = num_small_sp == 32'h1; // @[BFS.scala 921:42]
  wire [31:0] vertices_per_sp = num_small_sp == 32'h1 ? {{12'd0}, io_graph_scale[19:0]} : 32'h80000; // @[BFS.scala 921:28]
  wire [33:0] _GEN_51 = {vertices_per_sp, 2'h0}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T = {{13'd0}, _GEN_51}; // @[BFS.scala 924:35]
  wire [46:0] _wb_bram_T_2 = _wb_bram_T + 47'h4000; // @[BFS.scala 924:57]
  wire [31:0] _GEN_52 = {{12'd0}, io_graph_scale[19:0]}; // @[BFS.scala 926:36]
  wire [31:0] _wb_bram_T_5 = vertices_per_sp + _GEN_52; // @[BFS.scala 926:36]
  wire [33:0] _GEN_53 = {_wb_bram_T_5, 2'h0}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_6 = {{13'd0}, _GEN_53}; // @[BFS.scala 926:60]
  wire [46:0] _wb_bram_T_8 = _wb_bram_T_6 + 47'h4000; // @[BFS.scala 926:82]
  wire [34:0] _GEN_54 = {vertices_per_sp, 3'h0}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_9 = {{12'd0}, _GEN_54}; // @[BFS.scala 929:35]
  wire [46:0] _wb_bram_T_11 = _wb_bram_T_9 + 47'h4000; // @[BFS.scala 929:57]
  wire [46:0] _GEN_8 = num_small_sp == 32'h2 ? _wb_bram_T_8 : _wb_bram_T_11; // @[BFS.scala 925:37 BFS.scala 926:15 BFS.scala 929:15]
  wire [46:0] _GEN_9 = _vertices_per_sp_T ? _wb_bram_T_2 : _GEN_8; // @[BFS.scala 923:31 BFS.scala 924:15]
  wire [31:0] _wb_bram_T_14 = wb_bram - 32'h40; // @[BFS.scala 932:44]
  wire [31:0] _wb_bram_T_15 = wb_bram > 32'h40 ? _wb_bram_T_14 : 32'h0; // @[BFS.scala 932:19]
  wire [31:0] _GEN_10 = _T_7 ? _wb_bram_T_15 : wb_bram; // @[BFS.scala 931:28 BFS.scala 932:13 BFS.scala 910:24]
  wire [46:0] _GEN_11 = _T_10 & wb_bram == 32'h0 ? _GEN_9 : {{15'd0}, _GEN_10}; // @[BFS.scala 922:49]
  reg [31:0] ready_counter; // @[BFS.scala 936:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[BFS.scala 939:36]
  bitmap_0 bitmap_ ( // @[BFS.scala 802:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 803:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(arbi_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  Scatter_in_reg_slice scatter_in ( // @[BFS.scala 828:26]
    .aclk(scatter_in_aclk),
    .aresetn(scatter_in_aresetn),
    .s_axis_tdata(scatter_in_s_axis_tdata),
    .s_axis_tvalid(scatter_in_s_axis_tvalid),
    .s_axis_tkeep(scatter_in_s_axis_tkeep),
    .s_axis_tready(scatter_in_s_axis_tready),
    .s_axis_tlast(scatter_in_s_axis_tlast),
    .m_axis_tdata(scatter_in_m_axis_tdata),
    .m_axis_tvalid(scatter_in_m_axis_tvalid),
    .m_axis_tkeep(scatter_in_m_axis_tkeep),
    .m_axis_tready(scatter_in_m_axis_tready),
    .m_axis_tlast(scatter_in_m_axis_tlast)
  );
  vid_32_fifo vertex_in_fifo ( // @[BFS.scala 844:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  scatter_out_reg_slice vertex_out_fifo ( // @[BFS.scala 857:31]
    .aclk(vertex_out_fifo_aclk),
    .aresetn(vertex_out_fifo_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast)
  );
  assign io_xbar_in_ready = scatter_in_s_axis_tready; // @[BFS.scala 833:20]
  assign io_end = _T_9 & _vertices_per_sp_T; // @[BFS.scala 934:46]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 902:19]
  assign bitmap__clka = clock; // @[BFS.scala 900:33]
  assign bitmap__dina = bitmap_write_data_bits; // @[BFS.scala 901:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 898:17]
  assign bitmap__wea = bitmap_write_addr_valid & ~bitmap_write_addr_bits[31]; // @[BFS.scala 899:44]
  assign bitmap__addrb = _bitmap_io_addrb_T_14[16:0]; // @[BFS.scala 894:19]
  assign bitmap__clkb = clock; // @[BFS.scala 895:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 893:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = vertex_in_fifo_m_axis_tvalid; // @[BFS.scala 854:25]
  assign arbi_io_xbar_in_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign arbi_io_xbar_in_bits_tkeep = _arbi_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign arbi_io_xbar_in_bits_tlast = vertex_in_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign arbi_io_ddr_out_ready = ~halt; // @[BFS.scala 892:28]
  assign scatter_in_aclk = clock; // @[BFS.scala 829:37]
  assign scatter_in_aresetn = ~reset; // @[BFS.scala 830:28]
  assign scatter_in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign scatter_in_s_axis_tvalid = io_xbar_in_valid; // @[BFS.scala 832:31]
  assign scatter_in_s_axis_tkeep = {{48'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign scatter_in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign scatter_in_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[BFS.scala 851:31]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[BFS.scala 845:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 846:39]
  assign vertex_in_fifo_s_axis_tdata = scatter_in_m_axis_tdata; // @[BFS.scala 847:34]
  assign vertex_in_fifo_s_axis_tvalid = scatter_in_m_axis_tvalid & (filtered_keep_0 | filtered_keep_1 | filtered_keep_2
     | filtered_keep_3 | filtered_keep_4 | filtered_keep_5 | filtered_keep_6 | filtered_keep_7 | filtered_keep_8 |
    filtered_keep_9 | filtered_keep_10 | filtered_keep_11 | filtered_keep_12 | filtered_keep_13 | filtered_keep_14 |
    filtered_keep_15); // @[BFS.scala 849:66]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[BFS.scala 850:57]
  assign vertex_in_fifo_s_axis_tlast = scatter_in_m_axis_tlast; // @[BFS.scala 848:34]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = arbi_io_xbar_in_ready; // @[BFS.scala 855:35]
  assign vertex_out_fifo_aclk = clock; // @[BFS.scala 858:42]
  assign vertex_out_fifo_aresetn = ~reset; // @[BFS.scala 859:33]
  assign vertex_out_fifo_s_axis_tdata = bitmap_write_addr_bits; // @[BFS.scala 897:35]
  assign vertex_out_fifo_s_axis_tvalid = bitmap_write_addr_valid; // @[BFS.scala 896:36]
  assign vertex_out_fifo_s_axis_tkeep = 4'h0;
  assign vertex_out_fifo_s_axis_tlast = 1'h0;
  assign vertex_out_fifo_m_axis_tready = 1'h1; // @[BFS.scala 903:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 804:30]
      local_fpga_id <= 3'h0; // @[BFS.scala 804:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[BFS.scala 805:17]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_valid <= 1'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_valid <= arbi_io_ddr_out_valid; // @[BFS.scala 866:23]
    end
    if (reset) begin // @[BFS.scala 864:28]
      bitmap_wait_bits <= 32'h0; // @[BFS.scala 864:28]
    end else if (~halt) begin // @[BFS.scala 865:14]
      bitmap_wait_bits <= arbi_io_ddr_out_bits_tdata; // @[BFS.scala 867:22]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_valid <= 1'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_valid <= bitmap_wait_valid & _bitmap_write_addr_valid_T_9; // @[BFS.scala 872:29]
    end
    if (reset) begin // @[BFS.scala 870:34]
      bitmap_write_addr_bits <= 32'h0; // @[BFS.scala 870:34]
    end else if (_T) begin // @[BFS.scala 871:15]
      bitmap_write_addr_bits <= bitmap_wait_bits; // @[BFS.scala 874:28]
    end
    if (reset) begin // @[BFS.scala 876:34]
      bitmap_write_data_bits <= 9'h0; // @[BFS.scala 876:34]
    end else begin
      bitmap_write_data_bits <= _GEN_5[8:0];
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_valid <= 1'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_valid <= bitmap_write_addr_valid & arbi_io_ddr_out_valid &
        _bitmap_write_data_forward_valid_T_15; // @[BFS.scala 883:35]
    end
    if (reset) begin // @[BFS.scala 882:42]
      bitmap_write_data_forward_bits <= 9'h0; // @[BFS.scala 882:42]
    end else begin
      bitmap_write_data_forward_bits <= bitmap_write_data_bits; // @[BFS.scala 885:34]
    end
    if (reset) begin // @[BFS.scala 910:24]
      wb_bram <= 32'h0; // @[BFS.scala 910:24]
    end else begin
      wb_bram <= _GEN_11[31:0];
    end
    if (reset) begin // @[BFS.scala 914:29]
      num_small_sp <= 32'h0; // @[BFS.scala 914:29]
    end else if (vertex_out_fifo_m_axis_tvalid & vertex_out_fifo_m_axis_tdata[31]) begin // @[BFS.scala 915:96]
      num_small_sp <= _num_small_sp_T_3; // @[BFS.scala 916:18]
    end else if (wb_bram > 32'h0 & wb_bram <= 32'h40 & num_small_sp != 32'h0) begin // @[BFS.scala 918:71]
      num_small_sp <= _num_small_sp_T_5; // @[BFS.scala 919:18]
    end
    if (reset) begin // @[BFS.scala 936:30]
      ready_counter <= 32'h0; // @[BFS.scala 936:30]
    end else if (~io_xbar_in_ready & io_xbar_in_valid) begin // @[BFS.scala 938:68]
      ready_counter <= _ready_counter_T_1; // @[BFS.scala 939:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bitmap_wait_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bitmap_wait_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bitmap_write_addr_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bitmap_write_addr_bits = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bitmap_write_data_bits = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  bitmap_write_data_forward_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bitmap_write_data_forward_bits = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  wb_bram = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  num_small_sp = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ready_counter = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_arbitrator_16(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [127:0] io_xbar_in_bits_tdata,
  input  [3:0]   io_xbar_in_bits_tkeep,
  input          io_xbar_in_bits_tlast,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  in_aclk; // @[util.scala 455:18]
  wire  in_aresetn; // @[util.scala 455:18]
  wire [127:0] in_s_axis_tdata; // @[util.scala 455:18]
  wire  in_s_axis_tvalid; // @[util.scala 455:18]
  wire [15:0] in_s_axis_tkeep; // @[util.scala 455:18]
  wire  in_s_axis_tready; // @[util.scala 455:18]
  wire  in_s_axis_tlast; // @[util.scala 455:18]
  wire [127:0] in_m_axis_tdata; // @[util.scala 455:18]
  wire  in_m_axis_tvalid; // @[util.scala 455:18]
  wire [15:0] in_m_axis_tkeep; // @[util.scala 455:18]
  wire  in_m_axis_tready; // @[util.scala 455:18]
  wire  in_m_axis_tlast; // @[util.scala 455:18]
  wire  mid_aclk; // @[util.scala 465:19]
  wire  mid_aresetn; // @[util.scala 465:19]
  wire [127:0] mid_s_axis_tdata; // @[util.scala 465:19]
  wire  mid_s_axis_tvalid; // @[util.scala 465:19]
  wire [15:0] mid_s_axis_tkeep; // @[util.scala 465:19]
  wire  mid_s_axis_tready; // @[util.scala 465:19]
  wire  mid_s_axis_tlast; // @[util.scala 465:19]
  wire [127:0] mid_m_axis_tdata; // @[util.scala 465:19]
  wire  mid_m_axis_tvalid; // @[util.scala 465:19]
  wire [15:0] mid_m_axis_tkeep; // @[util.scala 465:19]
  wire  mid_m_axis_tready; // @[util.scala 465:19]
  wire  mid_m_axis_tlast; // @[util.scala 465:19]
  wire  out_aclk; // @[util.scala 485:19]
  wire  out_aresetn; // @[util.scala 485:19]
  wire [31:0] out_s_axis_tdata; // @[util.scala 485:19]
  wire  out_s_axis_tvalid; // @[util.scala 485:19]
  wire [3:0] out_s_axis_tkeep; // @[util.scala 485:19]
  wire  out_s_axis_tready; // @[util.scala 485:19]
  wire  out_s_axis_tlast; // @[util.scala 485:19]
  wire [31:0] out_m_axis_tdata; // @[util.scala 485:19]
  wire  out_m_axis_tvalid; // @[util.scala 485:19]
  wire [3:0] out_m_axis_tkeep; // @[util.scala 485:19]
  wire  out_m_axis_tready; // @[util.scala 485:19]
  wire  out_m_axis_tlast; // @[util.scala 485:19]
  wire  in_keep_0 = in_m_axis_tkeep[0]; // @[util.scala 463:97]
  wire  in_keep_1 = in_m_axis_tkeep[1]; // @[util.scala 463:97]
  wire  in_keep_2 = in_m_axis_tkeep[2]; // @[util.scala 463:97]
  wire  in_keep_3 = in_m_axis_tkeep[3]; // @[util.scala 463:97]
  wire [2:0] _in_count_WIRE = {{2'd0}, in_keep_0}; // @[util.scala 464:43 util.scala 464:43]
  wire [2:0] _in_count_WIRE_1 = {{2'd0}, in_keep_1}; // @[util.scala 464:43 util.scala 464:43]
  wire [2:0] _in_count_T_1 = _in_count_WIRE + _in_count_WIRE_1; // @[util.scala 464:82]
  wire [2:0] _in_count_WIRE_2 = {{2'd0}, in_keep_2}; // @[util.scala 464:43 util.scala 464:43]
  wire [2:0] _in_count_T_3 = _in_count_T_1 + _in_count_WIRE_2; // @[util.scala 464:82]
  wire [2:0] _in_count_WIRE_3 = {{2'd0}, in_keep_3}; // @[util.scala 464:43 util.scala 464:43]
  wire [2:0] in_count = _in_count_T_3 + _in_count_WIRE_3; // @[util.scala 464:82]
  wire [12:0] mid_io_s_axis_tkeep_lo = in_m_axis_tkeep[12:0]; // @[util.scala 472:58]
  wire  keep_0 = mid_m_axis_tkeep[0]; // @[util.scala 476:95]
  wire  keep_1 = mid_m_axis_tkeep[1]; // @[util.scala 476:95]
  wire  keep_2 = mid_m_axis_tkeep[2]; // @[util.scala 476:95]
  wire  keep_3 = mid_m_axis_tkeep[3]; // @[util.scala 476:95]
  reg  index_0; // @[util.scala 477:22]
  reg  index_1; // @[util.scala 477:22]
  reg  index_2; // @[util.scala 477:22]
  reg  index_3; // @[util.scala 477:22]
  wire  ungrant_keep_0 = keep_0 & ~index_0; // @[util.scala 479:22]
  wire  ungrant_keep_1 = keep_1 & ~index_1; // @[util.scala 479:22]
  wire  ungrant_keep_2 = keep_2 & ~index_2; // @[util.scala 479:22]
  wire  ungrant_keep_3 = keep_3 & ~index_3; // @[util.scala 479:22]
  wire  grant_1 = ~ungrant_keep_0; // @[util.scala 363:78]
  wire  grant_2 = ~(ungrant_keep_0 | ungrant_keep_1); // @[util.scala 363:78]
  wire  grant_3 = ~(ungrant_keep_0 | ungrant_keep_1 | ungrant_keep_2); // @[util.scala 363:78]
  wire  choosen_keep_1 = grant_1 & ungrant_keep_1; // @[util.scala 483:22]
  wire  choosen_keep_2 = grant_2 & ungrant_keep_2; // @[util.scala 483:22]
  wire  choosen_keep_3 = grant_3 & ungrant_keep_3; // @[util.scala 483:22]
  wire  _T_1 = mid_m_axis_tvalid; // @[util.scala 491:72]
  wire  _T_4 = out_s_axis_tready; // @[util.scala 493:78]
  wire  _T_5 = out_s_axis_tvalid & out_s_axis_tready; // @[util.scala 493:48]
  reg [2:0] count; // @[util.scala 499:22]
  wire [2:0] next_count = mid_m_axis_tkeep[15:13]; // @[util.scala 500:39]
  wire [2:0] _count_T_1 = next_count - 3'h1; // @[util.scala 503:27]
  wire [2:0] _count_T_3 = count - 3'h1; // @[util.scala 505:22]
  wire [31:0] _out_io_s_axis_tdata_T_4 = ungrant_keep_0 ? mid_m_axis_tdata[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_5 = choosen_keep_1 ? mid_m_axis_tdata[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_6 = choosen_keep_2 ? mid_m_axis_tdata[95:64] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_7 = choosen_keep_3 ? mid_m_axis_tdata[127:96] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_8 = _out_io_s_axis_tdata_T_4 | _out_io_s_axis_tdata_T_5; // @[Mux.scala 27:72]
  wire [31:0] _out_io_s_axis_tdata_T_9 = _out_io_s_axis_tdata_T_8 | _out_io_s_axis_tdata_T_6; // @[Mux.scala 27:72]
  axis_arbitrator_in_reg_slice_16 in ( // @[util.scala 455:18]
    .aclk(in_aclk),
    .aresetn(in_aresetn),
    .s_axis_tdata(in_s_axis_tdata),
    .s_axis_tvalid(in_s_axis_tvalid),
    .s_axis_tkeep(in_s_axis_tkeep),
    .s_axis_tready(in_s_axis_tready),
    .s_axis_tlast(in_s_axis_tlast),
    .m_axis_tdata(in_m_axis_tdata),
    .m_axis_tvalid(in_m_axis_tvalid),
    .m_axis_tkeep(in_m_axis_tkeep),
    .m_axis_tready(in_m_axis_tready),
    .m_axis_tlast(in_m_axis_tlast)
  );
  axis_arbitrator_in_reg_slice_16 mid ( // @[util.scala 465:19]
    .aclk(mid_aclk),
    .aresetn(mid_aresetn),
    .s_axis_tdata(mid_s_axis_tdata),
    .s_axis_tvalid(mid_s_axis_tvalid),
    .s_axis_tkeep(mid_s_axis_tkeep),
    .s_axis_tready(mid_s_axis_tready),
    .s_axis_tlast(mid_s_axis_tlast),
    .m_axis_tdata(mid_m_axis_tdata),
    .m_axis_tvalid(mid_m_axis_tvalid),
    .m_axis_tkeep(mid_m_axis_tkeep),
    .m_axis_tready(mid_m_axis_tready),
    .m_axis_tlast(mid_m_axis_tlast)
  );
  axis_arbitrator_out_reg_slice_4 out ( // @[util.scala 485:19]
    .aclk(out_aclk),
    .aresetn(out_aresetn),
    .s_axis_tdata(out_s_axis_tdata),
    .s_axis_tvalid(out_s_axis_tvalid),
    .s_axis_tkeep(out_s_axis_tkeep),
    .s_axis_tready(out_s_axis_tready),
    .s_axis_tlast(out_s_axis_tlast),
    .m_axis_tdata(out_m_axis_tdata),
    .m_axis_tvalid(out_m_axis_tvalid),
    .m_axis_tkeep(out_m_axis_tkeep),
    .m_axis_tready(out_m_axis_tready),
    .m_axis_tlast(out_m_axis_tlast)
  );
  assign io_xbar_in_ready = in_s_axis_tready; // @[util.scala 461:20]
  assign io_ddr_out_valid = out_m_axis_tvalid; // @[util.scala 516:20]
  assign io_ddr_out_bits_tdata = out_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign in_aclk = clock; // @[util.scala 457:29]
  assign in_aresetn = ~reset; // @[util.scala 458:20]
  assign in_s_axis_tdata = io_xbar_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_s_axis_tvalid = io_xbar_in_valid; // @[util.scala 460:23]
  assign in_s_axis_tkeep = {{12'd0}, io_xbar_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign in_s_axis_tlast = io_xbar_in_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign in_m_axis_tready = mid_s_axis_tready; // @[util.scala 473:23]
  assign mid_aclk = clock; // @[util.scala 467:30]
  assign mid_aresetn = ~reset; // @[util.scala 468:21]
  assign mid_s_axis_tdata = in_m_axis_tdata; // @[util.scala 470:23]
  assign mid_s_axis_tvalid = in_m_axis_tvalid; // @[util.scala 469:24]
  assign mid_s_axis_tkeep = {in_count,mid_io_s_axis_tkeep_lo}; // @[Cat.scala 30:58]
  assign mid_s_axis_tlast = in_m_axis_tlast; // @[util.scala 471:23]
  assign mid_m_axis_tready = _T_4 & (count == 3'h1 | next_count == 3'h1); // @[util.scala 508:57]
  assign out_aclk = clock; // @[util.scala 486:30]
  assign out_aresetn = ~reset; // @[util.scala 487:21]
  assign out_s_axis_tdata = _out_io_s_axis_tdata_T_9 | _out_io_s_axis_tdata_T_7; // @[Mux.scala 27:72]
  assign out_s_axis_tvalid = (ungrant_keep_0 | choosen_keep_1 | choosen_keep_2 | choosen_keep_3) & _T_1; // @[util.scala 510:52]
  assign out_s_axis_tkeep = 4'h1; // @[util.scala 511:23]
  assign out_s_axis_tlast = 1'h1; // @[util.scala 512:23]
  assign out_m_axis_tready = io_ddr_out_ready; // @[util.scala 517:24]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 477:22]
      index_0 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_0 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_0 <= index_0 | ungrant_keep_0; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_1 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_1 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_1 <= index_1 | choosen_keep_1; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_2 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_2 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_2 <= index_2 | choosen_keep_2; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 477:22]
      index_3 <= 1'h0; // @[util.scala 477:22]
    end else if (mid_m_axis_tready & mid_m_axis_tvalid) begin // @[util.scala 491:75]
      index_3 <= 1'h0; // @[util.scala 492:11]
    end else if (out_s_axis_tvalid & out_s_axis_tready) begin // @[util.scala 493:81]
      index_3 <= index_3 | choosen_keep_3; // @[util.scala 494:11]
    end
    if (reset) begin // @[util.scala 499:22]
      count <= 3'h0; // @[util.scala 499:22]
    end else if (_T_5) begin // @[util.scala 501:71]
      if (count == 3'h0) begin // @[util.scala 502:24]
        count <= _count_T_1; // @[util.scala 503:13]
      end else begin
        count <= _count_T_3; // @[util.scala 505:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  index_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  index_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  index_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  index_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  count = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Gather(
  input          clock,
  input          reset,
  output         io_ddr_in_ready,
  input          io_ddr_in_valid,
  input  [511:0] io_ddr_in_bits_tdata,
  input  [15:0]  io_ddr_in_bits_tkeep,
  input          io_gather_out_0_ready,
  output         io_gather_out_0_valid,
  output [31:0]  io_gather_out_0_bits_tdata,
  input          io_gather_out_1_ready,
  output         io_gather_out_1_valid,
  output [31:0]  io_gather_out_1_bits_tdata,
  input          io_gather_out_2_ready,
  output         io_gather_out_2_valid,
  output [31:0]  io_gather_out_2_bits_tdata,
  input          io_gather_out_3_ready,
  output         io_gather_out_3_valid,
  output [31:0]  io_gather_out_3_bits_tdata
);
  wire  broadcaster_aclk; // @[BFS.scala 205:27]
  wire  broadcaster_aresetn; // @[BFS.scala 205:27]
  wire [511:0] broadcaster_s_axis_tdata; // @[BFS.scala 205:27]
  wire  broadcaster_s_axis_tvalid; // @[BFS.scala 205:27]
  wire [63:0] broadcaster_s_axis_tkeep; // @[BFS.scala 205:27]
  wire  broadcaster_s_axis_tready; // @[BFS.scala 205:27]
  wire  broadcaster_s_axis_tlast; // @[BFS.scala 205:27]
  wire  broadcaster_s_axis_tid; // @[BFS.scala 205:27]
  wire [2559:0] broadcaster_m_axis_tdata; // @[BFS.scala 205:27]
  wire [4:0] broadcaster_m_axis_tvalid; // @[BFS.scala 205:27]
  wire [319:0] broadcaster_m_axis_tkeep; // @[BFS.scala 205:27]
  wire [4:0] broadcaster_m_axis_tready; // @[BFS.scala 205:27]
  wire [4:0] broadcaster_m_axis_tlast; // @[BFS.scala 205:27]
  wire [4:0] broadcaster_m_axis_tid; // @[BFS.scala 205:27]
  wire  v2Apply_fifo_aclk; // @[BFS.scala 212:28]
  wire  v2Apply_fifo_aresetn; // @[BFS.scala 212:28]
  wire [511:0] v2Apply_fifo_s_axis_tdata; // @[BFS.scala 212:28]
  wire  v2Apply_fifo_s_axis_tvalid; // @[BFS.scala 212:28]
  wire [63:0] v2Apply_fifo_s_axis_tkeep; // @[BFS.scala 212:28]
  wire  v2Apply_fifo_s_axis_tready; // @[BFS.scala 212:28]
  wire  v2Apply_fifo_s_axis_tlast; // @[BFS.scala 212:28]
  wire [511:0] v2Apply_fifo_m_axis_tdata; // @[BFS.scala 212:28]
  wire  v2Apply_fifo_m_axis_tvalid; // @[BFS.scala 212:28]
  wire [63:0] v2Apply_fifo_m_axis_tkeep; // @[BFS.scala 212:28]
  wire  v2Apply_fifo_m_axis_tready; // @[BFS.scala 212:28]
  wire  v2Apply_fifo_m_axis_tlast; // @[BFS.scala 212:28]
  wire  v2Broadcast_fifo_0_aclk; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_0_aresetn; // @[BFS.scala 221:16]
  wire [127:0] v2Broadcast_fifo_0_s_axis_tdata; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_0_s_axis_tvalid; // @[BFS.scala 221:16]
  wire [15:0] v2Broadcast_fifo_0_s_axis_tkeep; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_0_s_axis_tready; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_0_s_axis_tlast; // @[BFS.scala 221:16]
  wire [127:0] v2Broadcast_fifo_0_m_axis_tdata; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_0_m_axis_tvalid; // @[BFS.scala 221:16]
  wire [15:0] v2Broadcast_fifo_0_m_axis_tkeep; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_0_m_axis_tready; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_0_m_axis_tlast; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_1_aclk; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_1_aresetn; // @[BFS.scala 221:16]
  wire [127:0] v2Broadcast_fifo_1_s_axis_tdata; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_1_s_axis_tvalid; // @[BFS.scala 221:16]
  wire [15:0] v2Broadcast_fifo_1_s_axis_tkeep; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_1_s_axis_tready; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_1_s_axis_tlast; // @[BFS.scala 221:16]
  wire [127:0] v2Broadcast_fifo_1_m_axis_tdata; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_1_m_axis_tvalid; // @[BFS.scala 221:16]
  wire [15:0] v2Broadcast_fifo_1_m_axis_tkeep; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_1_m_axis_tready; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_1_m_axis_tlast; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_2_aclk; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_2_aresetn; // @[BFS.scala 221:16]
  wire [127:0] v2Broadcast_fifo_2_s_axis_tdata; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_2_s_axis_tvalid; // @[BFS.scala 221:16]
  wire [15:0] v2Broadcast_fifo_2_s_axis_tkeep; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_2_s_axis_tready; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_2_s_axis_tlast; // @[BFS.scala 221:16]
  wire [127:0] v2Broadcast_fifo_2_m_axis_tdata; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_2_m_axis_tvalid; // @[BFS.scala 221:16]
  wire [15:0] v2Broadcast_fifo_2_m_axis_tkeep; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_2_m_axis_tready; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_2_m_axis_tlast; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_3_aclk; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_3_aresetn; // @[BFS.scala 221:16]
  wire [127:0] v2Broadcast_fifo_3_s_axis_tdata; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_3_s_axis_tvalid; // @[BFS.scala 221:16]
  wire [15:0] v2Broadcast_fifo_3_s_axis_tkeep; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_3_s_axis_tready; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_3_s_axis_tlast; // @[BFS.scala 221:16]
  wire [127:0] v2Broadcast_fifo_3_m_axis_tdata; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_3_m_axis_tvalid; // @[BFS.scala 221:16]
  wire [15:0] v2Broadcast_fifo_3_m_axis_tkeep; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_3_m_axis_tready; // @[BFS.scala 221:16]
  wire  v2Broadcast_fifo_3_m_axis_tlast; // @[BFS.scala 221:16]
  wire  v2Broadcast_selecter_0_clock; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_0_reset; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_ready; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_valid; // @[BFS.scala 255:16]
  wire [127:0] v2Broadcast_selecter_0_io_xbar_in_bits_tdata; // @[BFS.scala 255:16]
  wire [3:0] v2Broadcast_selecter_0_io_xbar_in_bits_tkeep; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_bits_tlast; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_0_io_ddr_out_ready; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_0_io_ddr_out_valid; // @[BFS.scala 255:16]
  wire [31:0] v2Broadcast_selecter_0_io_ddr_out_bits_tdata; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_1_clock; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_1_reset; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_ready; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_valid; // @[BFS.scala 255:16]
  wire [127:0] v2Broadcast_selecter_1_io_xbar_in_bits_tdata; // @[BFS.scala 255:16]
  wire [3:0] v2Broadcast_selecter_1_io_xbar_in_bits_tkeep; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_bits_tlast; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_1_io_ddr_out_ready; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_1_io_ddr_out_valid; // @[BFS.scala 255:16]
  wire [31:0] v2Broadcast_selecter_1_io_ddr_out_bits_tdata; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_2_clock; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_2_reset; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_ready; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_valid; // @[BFS.scala 255:16]
  wire [127:0] v2Broadcast_selecter_2_io_xbar_in_bits_tdata; // @[BFS.scala 255:16]
  wire [3:0] v2Broadcast_selecter_2_io_xbar_in_bits_tkeep; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_bits_tlast; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_2_io_ddr_out_ready; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_2_io_ddr_out_valid; // @[BFS.scala 255:16]
  wire [31:0] v2Broadcast_selecter_2_io_ddr_out_bits_tdata; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_3_clock; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_3_reset; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_ready; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_valid; // @[BFS.scala 255:16]
  wire [127:0] v2Broadcast_selecter_3_io_xbar_in_bits_tdata; // @[BFS.scala 255:16]
  wire [3:0] v2Broadcast_selecter_3_io_xbar_in_bits_tkeep; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_bits_tlast; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_3_io_ddr_out_ready; // @[BFS.scala 255:16]
  wire  v2Broadcast_selecter_3_io_ddr_out_valid; // @[BFS.scala 255:16]
  wire [31:0] v2Broadcast_selecter_3_io_ddr_out_bits_tdata; // @[BFS.scala 255:16]
  wire [63:0] v2Broadcast_fifo_0_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[159:128],broadcaster_m_axis_tdata[31:0]}
    ; // @[BFS.scala 230:16]
  wire [63:0] v2Broadcast_fifo_0_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[415:384],broadcaster_m_axis_tdata[287:
    256]}; // @[BFS.scala 230:16]
  wire  _v2Broadcast_fifo_0_io_s_axis_tvalid_T_29 = broadcaster_m_axis_tkeep[0] | broadcaster_m_axis_tkeep[4] |
    broadcaster_m_axis_tkeep[8] | broadcaster_m_axis_tkeep[12]; // @[BFS.scala 240:17]
  wire [3:0] _v2Broadcast_fifo_0_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[12],broadcaster_m_axis_tkeep[8],
    broadcaster_m_axis_tkeep[4],broadcaster_m_axis_tkeep[0]}; // @[BFS.scala 243:16]
  wire [63:0] v2Broadcast_fifo_1_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[703:672],broadcaster_m_axis_tdata[575:
    544]}; // @[BFS.scala 230:16]
  wire [63:0] v2Broadcast_fifo_1_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[959:928],broadcaster_m_axis_tdata[831:
    800]}; // @[BFS.scala 230:16]
  wire  _v2Broadcast_fifo_1_io_s_axis_tvalid_T_30 = broadcaster_m_axis_tkeep[1] | broadcaster_m_axis_tkeep[5] |
    broadcaster_m_axis_tkeep[9] | broadcaster_m_axis_tkeep[13]; // @[BFS.scala 240:17]
  wire [3:0] _v2Broadcast_fifo_1_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[13],broadcaster_m_axis_tkeep[9],
    broadcaster_m_axis_tkeep[5],broadcaster_m_axis_tkeep[1]}; // @[BFS.scala 243:16]
  wire [63:0] v2Broadcast_fifo_2_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[1247:1216],broadcaster_m_axis_tdata[1119
    :1088]}; // @[BFS.scala 230:16]
  wire [63:0] v2Broadcast_fifo_2_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[1503:1472],broadcaster_m_axis_tdata[1375
    :1344]}; // @[BFS.scala 230:16]
  wire  _v2Broadcast_fifo_2_io_s_axis_tvalid_T_31 = broadcaster_m_axis_tkeep[2] | broadcaster_m_axis_tkeep[6] |
    broadcaster_m_axis_tkeep[10] | broadcaster_m_axis_tkeep[14]; // @[BFS.scala 240:17]
  wire [3:0] _v2Broadcast_fifo_2_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[14],broadcaster_m_axis_tkeep[10],
    broadcaster_m_axis_tkeep[6],broadcaster_m_axis_tkeep[2]}; // @[BFS.scala 243:16]
  wire [63:0] v2Broadcast_fifo_3_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[1791:1760],broadcaster_m_axis_tdata[1663
    :1632]}; // @[BFS.scala 230:16]
  wire [63:0] v2Broadcast_fifo_3_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[2047:2016],broadcaster_m_axis_tdata[1919
    :1888]}; // @[BFS.scala 230:16]
  wire  _v2Broadcast_fifo_3_io_s_axis_tvalid_T_32 = broadcaster_m_axis_tkeep[3] | broadcaster_m_axis_tkeep[7] |
    broadcaster_m_axis_tkeep[11] | broadcaster_m_axis_tkeep[15]; // @[BFS.scala 240:17]
  wire [3:0] _v2Broadcast_fifo_3_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[15],broadcaster_m_axis_tkeep[11],
    broadcaster_m_axis_tkeep[7],broadcaster_m_axis_tkeep[3]}; // @[BFS.scala 243:16]
  wire  _broadcaster_io_m_axis_tready_WIRE_1 = v2Broadcast_fifo_1_s_axis_tready; // @[BFS.scala 248:101 BFS.scala 248:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_0 = v2Broadcast_fifo_0_s_axis_tready; // @[BFS.scala 248:101 BFS.scala 248:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_3 = v2Broadcast_fifo_3_s_axis_tready; // @[BFS.scala 248:101 BFS.scala 248:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_2 = v2Broadcast_fifo_2_s_axis_tready; // @[BFS.scala 248:101 BFS.scala 248:101]
  wire [3:0] broadcaster_io_m_axis_tready_lo_1 = {_broadcaster_io_m_axis_tready_WIRE_3,
    _broadcaster_io_m_axis_tready_WIRE_2,_broadcaster_io_m_axis_tready_WIRE_1,_broadcaster_io_m_axis_tready_WIRE_0}; // @[BFS.scala 248:151]
  wire [15:0] _v2Broadcast_selecter_0_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_0_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [15:0] _v2Broadcast_selecter_1_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_1_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [15:0] _v2Broadcast_selecter_2_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_2_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [15:0] _v2Broadcast_selecter_3_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_3_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  gather_broadcaster broadcaster ( // @[BFS.scala 205:27]
    .aclk(broadcaster_aclk),
    .aresetn(broadcaster_aresetn),
    .s_axis_tdata(broadcaster_s_axis_tdata),
    .s_axis_tvalid(broadcaster_s_axis_tvalid),
    .s_axis_tkeep(broadcaster_s_axis_tkeep),
    .s_axis_tready(broadcaster_s_axis_tready),
    .s_axis_tlast(broadcaster_s_axis_tlast),
    .s_axis_tid(broadcaster_s_axis_tid),
    .m_axis_tdata(broadcaster_m_axis_tdata),
    .m_axis_tvalid(broadcaster_m_axis_tvalid),
    .m_axis_tkeep(broadcaster_m_axis_tkeep),
    .m_axis_tready(broadcaster_m_axis_tready),
    .m_axis_tlast(broadcaster_m_axis_tlast),
    .m_axis_tid(broadcaster_m_axis_tid)
  );
  v2A_reg_slice v2Apply_fifo ( // @[BFS.scala 212:28]
    .aclk(v2Apply_fifo_aclk),
    .aresetn(v2Apply_fifo_aresetn),
    .s_axis_tdata(v2Apply_fifo_s_axis_tdata),
    .s_axis_tvalid(v2Apply_fifo_s_axis_tvalid),
    .s_axis_tkeep(v2Apply_fifo_s_axis_tkeep),
    .s_axis_tready(v2Apply_fifo_s_axis_tready),
    .s_axis_tlast(v2Apply_fifo_s_axis_tlast),
    .m_axis_tdata(v2Apply_fifo_m_axis_tdata),
    .m_axis_tvalid(v2Apply_fifo_m_axis_tvalid),
    .m_axis_tkeep(v2Apply_fifo_m_axis_tkeep),
    .m_axis_tready(v2Apply_fifo_m_axis_tready),
    .m_axis_tlast(v2Apply_fifo_m_axis_tlast)
  );
  v2B_reg_slice v2Broadcast_fifo_0 ( // @[BFS.scala 221:16]
    .aclk(v2Broadcast_fifo_0_aclk),
    .aresetn(v2Broadcast_fifo_0_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_0_s_axis_tdata),
    .s_axis_tvalid(v2Broadcast_fifo_0_s_axis_tvalid),
    .s_axis_tkeep(v2Broadcast_fifo_0_s_axis_tkeep),
    .s_axis_tready(v2Broadcast_fifo_0_s_axis_tready),
    .s_axis_tlast(v2Broadcast_fifo_0_s_axis_tlast),
    .m_axis_tdata(v2Broadcast_fifo_0_m_axis_tdata),
    .m_axis_tvalid(v2Broadcast_fifo_0_m_axis_tvalid),
    .m_axis_tkeep(v2Broadcast_fifo_0_m_axis_tkeep),
    .m_axis_tready(v2Broadcast_fifo_0_m_axis_tready),
    .m_axis_tlast(v2Broadcast_fifo_0_m_axis_tlast)
  );
  v2B_reg_slice v2Broadcast_fifo_1 ( // @[BFS.scala 221:16]
    .aclk(v2Broadcast_fifo_1_aclk),
    .aresetn(v2Broadcast_fifo_1_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_1_s_axis_tdata),
    .s_axis_tvalid(v2Broadcast_fifo_1_s_axis_tvalid),
    .s_axis_tkeep(v2Broadcast_fifo_1_s_axis_tkeep),
    .s_axis_tready(v2Broadcast_fifo_1_s_axis_tready),
    .s_axis_tlast(v2Broadcast_fifo_1_s_axis_tlast),
    .m_axis_tdata(v2Broadcast_fifo_1_m_axis_tdata),
    .m_axis_tvalid(v2Broadcast_fifo_1_m_axis_tvalid),
    .m_axis_tkeep(v2Broadcast_fifo_1_m_axis_tkeep),
    .m_axis_tready(v2Broadcast_fifo_1_m_axis_tready),
    .m_axis_tlast(v2Broadcast_fifo_1_m_axis_tlast)
  );
  v2B_reg_slice v2Broadcast_fifo_2 ( // @[BFS.scala 221:16]
    .aclk(v2Broadcast_fifo_2_aclk),
    .aresetn(v2Broadcast_fifo_2_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_2_s_axis_tdata),
    .s_axis_tvalid(v2Broadcast_fifo_2_s_axis_tvalid),
    .s_axis_tkeep(v2Broadcast_fifo_2_s_axis_tkeep),
    .s_axis_tready(v2Broadcast_fifo_2_s_axis_tready),
    .s_axis_tlast(v2Broadcast_fifo_2_s_axis_tlast),
    .m_axis_tdata(v2Broadcast_fifo_2_m_axis_tdata),
    .m_axis_tvalid(v2Broadcast_fifo_2_m_axis_tvalid),
    .m_axis_tkeep(v2Broadcast_fifo_2_m_axis_tkeep),
    .m_axis_tready(v2Broadcast_fifo_2_m_axis_tready),
    .m_axis_tlast(v2Broadcast_fifo_2_m_axis_tlast)
  );
  v2B_reg_slice v2Broadcast_fifo_3 ( // @[BFS.scala 221:16]
    .aclk(v2Broadcast_fifo_3_aclk),
    .aresetn(v2Broadcast_fifo_3_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_3_s_axis_tdata),
    .s_axis_tvalid(v2Broadcast_fifo_3_s_axis_tvalid),
    .s_axis_tkeep(v2Broadcast_fifo_3_s_axis_tkeep),
    .s_axis_tready(v2Broadcast_fifo_3_s_axis_tready),
    .s_axis_tlast(v2Broadcast_fifo_3_s_axis_tlast),
    .m_axis_tdata(v2Broadcast_fifo_3_m_axis_tdata),
    .m_axis_tvalid(v2Broadcast_fifo_3_m_axis_tvalid),
    .m_axis_tkeep(v2Broadcast_fifo_3_m_axis_tkeep),
    .m_axis_tready(v2Broadcast_fifo_3_m_axis_tready),
    .m_axis_tlast(v2Broadcast_fifo_3_m_axis_tlast)
  );
  axis_arbitrator_16 v2Broadcast_selecter_0 ( // @[BFS.scala 255:16]
    .clock(v2Broadcast_selecter_0_clock),
    .reset(v2Broadcast_selecter_0_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_0_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_0_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(v2Broadcast_selecter_0_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(v2Broadcast_selecter_0_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_0_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_0_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_16 v2Broadcast_selecter_1 ( // @[BFS.scala 255:16]
    .clock(v2Broadcast_selecter_1_clock),
    .reset(v2Broadcast_selecter_1_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_1_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_1_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(v2Broadcast_selecter_1_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(v2Broadcast_selecter_1_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_1_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_1_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_16 v2Broadcast_selecter_2 ( // @[BFS.scala 255:16]
    .clock(v2Broadcast_selecter_2_clock),
    .reset(v2Broadcast_selecter_2_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_2_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_2_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(v2Broadcast_selecter_2_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(v2Broadcast_selecter_2_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_2_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_2_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_16 v2Broadcast_selecter_3 ( // @[BFS.scala 255:16]
    .clock(v2Broadcast_selecter_3_clock),
    .reset(v2Broadcast_selecter_3_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_3_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_3_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(v2Broadcast_selecter_3_io_xbar_in_bits_tlast),
    .io_ddr_out_ready(v2Broadcast_selecter_3_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_3_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_3_io_ddr_out_bits_tdata)
  );
  assign io_ddr_in_ready = broadcaster_s_axis_tready; // @[BFS.scala 208:19]
  assign io_gather_out_0_valid = v2Broadcast_selecter_0_io_ddr_out_valid; // @[BFS.scala 262:20]
  assign io_gather_out_0_bits_tdata = v2Broadcast_selecter_0_io_ddr_out_bits_tdata; // @[BFS.scala 262:20]
  assign io_gather_out_1_valid = v2Broadcast_selecter_1_io_ddr_out_valid; // @[BFS.scala 262:20]
  assign io_gather_out_1_bits_tdata = v2Broadcast_selecter_1_io_ddr_out_bits_tdata; // @[BFS.scala 262:20]
  assign io_gather_out_2_valid = v2Broadcast_selecter_2_io_ddr_out_valid; // @[BFS.scala 262:20]
  assign io_gather_out_2_bits_tdata = v2Broadcast_selecter_2_io_ddr_out_bits_tdata; // @[BFS.scala 262:20]
  assign io_gather_out_3_valid = v2Broadcast_selecter_3_io_ddr_out_valid; // @[BFS.scala 262:20]
  assign io_gather_out_3_bits_tdata = v2Broadcast_selecter_3_io_ddr_out_bits_tdata; // @[BFS.scala 262:20]
  assign broadcaster_aclk = clock; // @[BFS.scala 210:38]
  assign broadcaster_aresetn = ~reset; // @[BFS.scala 209:29]
  assign broadcaster_s_axis_tdata = io_ddr_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign broadcaster_s_axis_tvalid = io_ddr_in_valid; // @[BFS.scala 207:32]
  assign broadcaster_s_axis_tkeep = {{48'd0}, io_ddr_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign broadcaster_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign broadcaster_s_axis_tid = 1'h0;
  assign broadcaster_m_axis_tready = {v2Apply_fifo_s_axis_tready,broadcaster_io_m_axis_tready_lo_1}; // @[Cat.scala 30:58]
  assign v2Apply_fifo_aclk = clock; // @[BFS.scala 213:39]
  assign v2Apply_fifo_aresetn = ~reset; // @[BFS.scala 214:30]
  assign v2Apply_fifo_s_axis_tdata = broadcaster_m_axis_tdata[2559:2048]; // @[BFS.scala 215:62]
  assign v2Apply_fifo_s_axis_tvalid = broadcaster_m_axis_tvalid[4]; // @[BFS.scala 216:64]
  assign v2Apply_fifo_s_axis_tkeep = broadcaster_m_axis_tkeep[319:256]; // @[BFS.scala 217:62]
  assign v2Apply_fifo_s_axis_tlast = broadcaster_m_axis_tlast[4]; // @[BFS.scala 218:62]
  assign v2Apply_fifo_m_axis_tready = 1'h1; // @[BFS.scala 251:33]
  assign v2Broadcast_fifo_0_aclk = clock; // @[BFS.scala 226:32]
  assign v2Broadcast_fifo_0_aresetn = ~reset; // @[BFS.scala 225:23]
  assign v2Broadcast_fifo_0_s_axis_tdata = {v2Broadcast_fifo_0_io_s_axis_tdata_hi,v2Broadcast_fifo_0_io_s_axis_tdata_lo}
    ; // @[BFS.scala 230:16]
  assign v2Broadcast_fifo_0_s_axis_tvalid = broadcaster_m_axis_tvalid[0] & _v2Broadcast_fifo_0_io_s_axis_tvalid_T_29; // @[BFS.scala 231:61]
  assign v2Broadcast_fifo_0_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_0_io_s_axis_tkeep_T_9}; // @[BFS.scala 243:16]
  assign v2Broadcast_fifo_0_s_axis_tlast = broadcaster_m_axis_tlast[0]; // @[BFS.scala 244:55]
  assign v2Broadcast_fifo_0_m_axis_tready = v2Broadcast_selecter_0_io_xbar_in_ready; // @[BFS.scala 261:44]
  assign v2Broadcast_fifo_1_aclk = clock; // @[BFS.scala 226:32]
  assign v2Broadcast_fifo_1_aresetn = ~reset; // @[BFS.scala 225:23]
  assign v2Broadcast_fifo_1_s_axis_tdata = {v2Broadcast_fifo_1_io_s_axis_tdata_hi,v2Broadcast_fifo_1_io_s_axis_tdata_lo}
    ; // @[BFS.scala 230:16]
  assign v2Broadcast_fifo_1_s_axis_tvalid = broadcaster_m_axis_tvalid[1] & _v2Broadcast_fifo_1_io_s_axis_tvalid_T_30; // @[BFS.scala 231:61]
  assign v2Broadcast_fifo_1_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_1_io_s_axis_tkeep_T_9}; // @[BFS.scala 243:16]
  assign v2Broadcast_fifo_1_s_axis_tlast = broadcaster_m_axis_tlast[1]; // @[BFS.scala 244:55]
  assign v2Broadcast_fifo_1_m_axis_tready = v2Broadcast_selecter_1_io_xbar_in_ready; // @[BFS.scala 261:44]
  assign v2Broadcast_fifo_2_aclk = clock; // @[BFS.scala 226:32]
  assign v2Broadcast_fifo_2_aresetn = ~reset; // @[BFS.scala 225:23]
  assign v2Broadcast_fifo_2_s_axis_tdata = {v2Broadcast_fifo_2_io_s_axis_tdata_hi,v2Broadcast_fifo_2_io_s_axis_tdata_lo}
    ; // @[BFS.scala 230:16]
  assign v2Broadcast_fifo_2_s_axis_tvalid = broadcaster_m_axis_tvalid[2] & _v2Broadcast_fifo_2_io_s_axis_tvalid_T_31; // @[BFS.scala 231:61]
  assign v2Broadcast_fifo_2_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_2_io_s_axis_tkeep_T_9}; // @[BFS.scala 243:16]
  assign v2Broadcast_fifo_2_s_axis_tlast = broadcaster_m_axis_tlast[2]; // @[BFS.scala 244:55]
  assign v2Broadcast_fifo_2_m_axis_tready = v2Broadcast_selecter_2_io_xbar_in_ready; // @[BFS.scala 261:44]
  assign v2Broadcast_fifo_3_aclk = clock; // @[BFS.scala 226:32]
  assign v2Broadcast_fifo_3_aresetn = ~reset; // @[BFS.scala 225:23]
  assign v2Broadcast_fifo_3_s_axis_tdata = {v2Broadcast_fifo_3_io_s_axis_tdata_hi,v2Broadcast_fifo_3_io_s_axis_tdata_lo}
    ; // @[BFS.scala 230:16]
  assign v2Broadcast_fifo_3_s_axis_tvalid = broadcaster_m_axis_tvalid[3] & _v2Broadcast_fifo_3_io_s_axis_tvalid_T_32; // @[BFS.scala 231:61]
  assign v2Broadcast_fifo_3_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_3_io_s_axis_tkeep_T_9}; // @[BFS.scala 243:16]
  assign v2Broadcast_fifo_3_s_axis_tlast = broadcaster_m_axis_tlast[3]; // @[BFS.scala 244:55]
  assign v2Broadcast_fifo_3_m_axis_tready = v2Broadcast_selecter_3_io_xbar_in_ready; // @[BFS.scala 261:44]
  assign v2Broadcast_selecter_0_clock = clock;
  assign v2Broadcast_selecter_0_reset = reset;
  assign v2Broadcast_selecter_0_io_xbar_in_valid = v2Broadcast_fifo_0_m_axis_tvalid; // @[BFS.scala 259:26]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tdata = v2Broadcast_fifo_0_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_0_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tlast = v2Broadcast_fifo_0_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign v2Broadcast_selecter_0_io_ddr_out_ready = io_gather_out_0_ready; // @[BFS.scala 262:20]
  assign v2Broadcast_selecter_1_clock = clock;
  assign v2Broadcast_selecter_1_reset = reset;
  assign v2Broadcast_selecter_1_io_xbar_in_valid = v2Broadcast_fifo_1_m_axis_tvalid; // @[BFS.scala 259:26]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tdata = v2Broadcast_fifo_1_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_1_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tlast = v2Broadcast_fifo_1_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign v2Broadcast_selecter_1_io_ddr_out_ready = io_gather_out_1_ready; // @[BFS.scala 262:20]
  assign v2Broadcast_selecter_2_clock = clock;
  assign v2Broadcast_selecter_2_reset = reset;
  assign v2Broadcast_selecter_2_io_xbar_in_valid = v2Broadcast_fifo_2_m_axis_tvalid; // @[BFS.scala 259:26]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tdata = v2Broadcast_fifo_2_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_2_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tlast = v2Broadcast_fifo_2_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign v2Broadcast_selecter_2_io_ddr_out_ready = io_gather_out_2_ready; // @[BFS.scala 262:20]
  assign v2Broadcast_selecter_3_clock = clock;
  assign v2Broadcast_selecter_3_reset = reset;
  assign v2Broadcast_selecter_3_io_xbar_in_valid = v2Broadcast_fifo_3_m_axis_tvalid; // @[BFS.scala 259:26]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tdata = v2Broadcast_fifo_3_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_3_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tlast = v2Broadcast_fifo_3_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign v2Broadcast_selecter_3_io_ddr_out_ready = io_gather_out_3_ready; // @[BFS.scala 262:20]
endmodule
module Apply(
  output  io_end,
  input   io_flush
);
  assign io_end = io_flush; // @[BFS.scala 196:10]
endmodule
module regFile(
  input         clock,
  input         reset,
  input  [63:0] io_dataIn,
  output [63:0] io_dataOut,
  input         io_writeFlag,
  input  [4:0]  io_rptr,
  input  [4:0]  io_wptr
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0; // @[util.scala 178:21]
  reg [63:0] regs_1; // @[util.scala 178:21]
  reg [63:0] regs_2; // @[util.scala 178:21]
  reg [63:0] regs_3; // @[util.scala 178:21]
  reg [63:0] regs_4; // @[util.scala 178:21]
  reg [63:0] regs_5; // @[util.scala 178:21]
  reg [63:0] regs_6; // @[util.scala 178:21]
  reg [63:0] regs_7; // @[util.scala 178:21]
  reg [63:0] regs_8; // @[util.scala 178:21]
  reg [63:0] regs_9; // @[util.scala 178:21]
  reg [63:0] regs_10; // @[util.scala 178:21]
  reg [63:0] regs_11; // @[util.scala 178:21]
  reg [63:0] regs_12; // @[util.scala 178:21]
  reg [63:0] regs_13; // @[util.scala 178:21]
  reg [63:0] regs_14; // @[util.scala 178:21]
  reg [63:0] regs_15; // @[util.scala 178:21]
  reg [63:0] regs_16; // @[util.scala 178:21]
  reg [63:0] regs_17; // @[util.scala 178:21]
  reg [63:0] regs_18; // @[util.scala 178:21]
  reg [63:0] regs_19; // @[util.scala 178:21]
  reg [63:0] regs_20; // @[util.scala 178:21]
  reg [63:0] regs_21; // @[util.scala 178:21]
  reg [63:0] regs_22; // @[util.scala 178:21]
  reg [63:0] regs_23; // @[util.scala 178:21]
  reg [63:0] regs_24; // @[util.scala 178:21]
  reg [63:0] regs_25; // @[util.scala 178:21]
  reg [63:0] regs_26; // @[util.scala 178:21]
  reg [63:0] regs_27; // @[util.scala 178:21]
  reg [63:0] regs_28; // @[util.scala 178:21]
  reg [63:0] regs_29; // @[util.scala 178:21]
  reg [63:0] regs_30; // @[util.scala 178:21]
  reg [63:0] regs_31; // @[util.scala 178:21]
  wire [63:0] _GEN_1 = 5'h1 == io_rptr ? regs_1 : regs_0; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_2 = 5'h2 == io_rptr ? regs_2 : _GEN_1; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_3 = 5'h3 == io_rptr ? regs_3 : _GEN_2; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_4 = 5'h4 == io_rptr ? regs_4 : _GEN_3; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_5 = 5'h5 == io_rptr ? regs_5 : _GEN_4; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_6 = 5'h6 == io_rptr ? regs_6 : _GEN_5; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_7 = 5'h7 == io_rptr ? regs_7 : _GEN_6; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_8 = 5'h8 == io_rptr ? regs_8 : _GEN_7; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_9 = 5'h9 == io_rptr ? regs_9 : _GEN_8; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_10 = 5'ha == io_rptr ? regs_10 : _GEN_9; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_11 = 5'hb == io_rptr ? regs_11 : _GEN_10; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_12 = 5'hc == io_rptr ? regs_12 : _GEN_11; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_13 = 5'hd == io_rptr ? regs_13 : _GEN_12; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_14 = 5'he == io_rptr ? regs_14 : _GEN_13; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_15 = 5'hf == io_rptr ? regs_15 : _GEN_14; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_16 = 5'h10 == io_rptr ? regs_16 : _GEN_15; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_17 = 5'h11 == io_rptr ? regs_17 : _GEN_16; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_18 = 5'h12 == io_rptr ? regs_18 : _GEN_17; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_19 = 5'h13 == io_rptr ? regs_19 : _GEN_18; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_20 = 5'h14 == io_rptr ? regs_20 : _GEN_19; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_21 = 5'h15 == io_rptr ? regs_21 : _GEN_20; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_22 = 5'h16 == io_rptr ? regs_22 : _GEN_21; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_23 = 5'h17 == io_rptr ? regs_23 : _GEN_22; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_24 = 5'h18 == io_rptr ? regs_24 : _GEN_23; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_25 = 5'h19 == io_rptr ? regs_25 : _GEN_24; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_26 = 5'h1a == io_rptr ? regs_26 : _GEN_25; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_27 = 5'h1b == io_rptr ? regs_27 : _GEN_26; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_28 = 5'h1c == io_rptr ? regs_28 : _GEN_27; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_29 = 5'h1d == io_rptr ? regs_29 : _GEN_28; // @[util.scala 180:14 util.scala 180:14]
  wire [63:0] _GEN_30 = 5'h1e == io_rptr ? regs_30 : _GEN_29; // @[util.scala 180:14 util.scala 180:14]
  assign io_dataOut = 5'h1f == io_rptr ? regs_31 : _GEN_30; // @[util.scala 180:14 util.scala 180:14]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 178:21]
      regs_0 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h0 == io_wptr) begin // @[util.scala 183:19]
        regs_0 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_1 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1 == io_wptr) begin // @[util.scala 183:19]
        regs_1 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_2 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h2 == io_wptr) begin // @[util.scala 183:19]
        regs_2 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_3 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h3 == io_wptr) begin // @[util.scala 183:19]
        regs_3 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_4 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h4 == io_wptr) begin // @[util.scala 183:19]
        regs_4 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_5 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h5 == io_wptr) begin // @[util.scala 183:19]
        regs_5 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_6 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h6 == io_wptr) begin // @[util.scala 183:19]
        regs_6 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_7 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h7 == io_wptr) begin // @[util.scala 183:19]
        regs_7 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_8 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h8 == io_wptr) begin // @[util.scala 183:19]
        regs_8 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_9 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h9 == io_wptr) begin // @[util.scala 183:19]
        regs_9 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_10 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'ha == io_wptr) begin // @[util.scala 183:19]
        regs_10 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_11 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hb == io_wptr) begin // @[util.scala 183:19]
        regs_11 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_12 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hc == io_wptr) begin // @[util.scala 183:19]
        regs_12 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_13 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hd == io_wptr) begin // @[util.scala 183:19]
        regs_13 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_14 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'he == io_wptr) begin // @[util.scala 183:19]
        regs_14 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_15 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hf == io_wptr) begin // @[util.scala 183:19]
        regs_15 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_16 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h10 == io_wptr) begin // @[util.scala 183:19]
        regs_16 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_17 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h11 == io_wptr) begin // @[util.scala 183:19]
        regs_17 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_18 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h12 == io_wptr) begin // @[util.scala 183:19]
        regs_18 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_19 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h13 == io_wptr) begin // @[util.scala 183:19]
        regs_19 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_20 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h14 == io_wptr) begin // @[util.scala 183:19]
        regs_20 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_21 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h15 == io_wptr) begin // @[util.scala 183:19]
        regs_21 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_22 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h16 == io_wptr) begin // @[util.scala 183:19]
        regs_22 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_23 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h17 == io_wptr) begin // @[util.scala 183:19]
        regs_23 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_24 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h18 == io_wptr) begin // @[util.scala 183:19]
        regs_24 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_25 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h19 == io_wptr) begin // @[util.scala 183:19]
        regs_25 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_26 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1a == io_wptr) begin // @[util.scala 183:19]
        regs_26 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_27 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1b == io_wptr) begin // @[util.scala 183:19]
        regs_27 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_28 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1c == io_wptr) begin // @[util.scala 183:19]
        regs_28 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_29 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1d == io_wptr) begin // @[util.scala 183:19]
        regs_29 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_30 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1e == io_wptr) begin // @[util.scala 183:19]
        regs_30 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_31 <= 64'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1f == io_wptr) begin // @[util.scala 183:19]
        regs_31 <= io_dataIn; // @[util.scala 183:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regs_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regs_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regs_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regs_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regs_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regs_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regs_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regs_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regs_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regs_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regs_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regs_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regs_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regs_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regs_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regs_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regs_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regs_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regs_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regs_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regs_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regs_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regs_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regs_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regs_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regs_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regs_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regs_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regs_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regs_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module readEdge_engine(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_rdata,
  input  [5:0]   io_in_bits_rid,
  input          io_in_bits_rlast,
  input          io_out_ready,
  output         io_out_valid,
  output [63:0]  io_out_bits_araddr,
  output [5:0]   io_out_bits_arid,
  output [7:0]   io_out_bits_arlen,
  output [2:0]   io_out_bits_arsize,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_edge_base_addr,
  output         io_read_edge_fifo_empty,
  output [7:0]   io_credit,
  input          io_credit_dec,
  output [63:0]  io_traveled_edges,
  input          io_signal
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  num_regfile_clock; // @[BFS.scala 341:27]
  wire  num_regfile_reset; // @[BFS.scala 341:27]
  wire [63:0] num_regfile_io_dataIn; // @[BFS.scala 341:27]
  wire [63:0] num_regfile_io_dataOut; // @[BFS.scala 341:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 341:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 341:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 341:27]
  wire  edge_read_buffer__full; // @[BFS.scala 387:32]
  wire [71:0] edge_read_buffer__din; // @[BFS.scala 387:32]
  wire  edge_read_buffer__wr_en; // @[BFS.scala 387:32]
  wire  edge_read_buffer__empty; // @[BFS.scala 387:32]
  wire [71:0] edge_read_buffer__dout; // @[BFS.scala 387:32]
  wire  edge_read_buffer__rd_en; // @[BFS.scala 387:32]
  wire [5:0] edge_read_buffer__data_count; // @[BFS.scala 387:32]
  wire  edge_read_buffer__clk; // @[BFS.scala 387:32]
  wire  edge_read_buffer__srst; // @[BFS.scala 387:32]
  wire  edge_read_buffer__valid; // @[BFS.scala 387:32]
  wire  free_queue_full; // @[BFS.scala 437:26]
  wire [5:0] free_queue_din; // @[BFS.scala 437:26]
  wire  free_queue_wr_en; // @[BFS.scala 437:26]
  wire  free_queue_empty; // @[BFS.scala 437:26]
  wire [5:0] free_queue_dout; // @[BFS.scala 437:26]
  wire  free_queue_rd_en; // @[BFS.scala 437:26]
  wire [5:0] free_queue_data_count; // @[BFS.scala 437:26]
  wire  free_queue_clk; // @[BFS.scala 437:26]
  wire  free_queue_srst; // @[BFS.scala 437:26]
  wire  free_queue_valid; // @[BFS.scala 437:26]
  reg [1:0] status; // @[BFS.scala 317:23]
  reg [31:0] num; // @[BFS.scala 318:20]
  wire  _T = status == 2'h0; // @[BFS.scala 319:15]
  wire  _T_2 = status == 2'h0 & io_in_valid & io_in_ready; // @[BFS.scala 319:48]
  wire  _T_6 = status == 2'h2; // @[BFS.scala 327:22]
  wire  _T_7 = status == 2'h1; // @[BFS.scala 327:60]
  wire  _T_8 = status == 2'h2 | status == 2'h1; // @[BFS.scala 327:50]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 331:35]
  wire  _T_13 = io_in_valid & io_in_ready; // @[BFS.scala 334:26]
  wire  _T_16 = ~io_in_bits_rid[5]; // @[BFS.scala 334:44]
  wire  _T_17 = io_in_valid & io_in_ready & ~io_in_bits_rid[5]; // @[BFS.scala 334:41]
  wire [63:0] _GEN_130 = {{32'd0}, io_in_bits_rdata[63:32]}; // @[BFS.scala 336:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_130; // @[BFS.scala 336:46]
  wire [31:0] _num_T_4 = num_regfile_io_dataOut[63:32] - 32'h4; // @[BFS.scala 345:103]
  wire [31:0] _num_T_10 = io_in_bits_rdata[63:32] - 32'h2; // @[BFS.scala 348:42]
  wire [31:0] _num_T_13 = num - 32'h4; // @[BFS.scala 354:18]
  wire [31:0] _num_T_17 = num > 32'h4 ? _num_T_13 : 32'h0; // @[BFS.scala 360:17]
  wire [31:0] _GEN_8 = io_in_bits_rlast ? 32'h0 : _num_T_17; // @[BFS.scala 357:36 BFS.scala 358:11 BFS.scala 360:11]
  wire  _GEN_12 = _T_8 & num > 32'h0; // @[BFS.scala 376:94 BFS.scala 377:11 BFS.scala 367:9]
  wire  _GEN_13 = _T & _T_16 ? 1'h0 : _GEN_12; // @[BFS.scala 370:72 BFS.scala 372:13]
  wire  keep_0 = _T & io_in_bits_rid[5] ? num_regfile_io_dataOut[63:32] > 32'h0 : _GEN_13; // @[BFS.scala 368:65 BFS.scala 369:11]
  wire  _GEN_15 = _T_8 & num > 32'h1; // @[BFS.scala 376:94 BFS.scala 377:11 BFS.scala 367:9]
  wire  _GEN_16 = _T & _T_16 ? 1'h0 : _GEN_15; // @[BFS.scala 370:72 BFS.scala 372:13]
  wire  keep_1 = _T & io_in_bits_rid[5] ? num_regfile_io_dataOut[63:32] > 32'h1 : _GEN_16; // @[BFS.scala 368:65 BFS.scala 369:11]
  wire  _GEN_18 = _T_8 & num > 32'h2; // @[BFS.scala 376:94 BFS.scala 377:11 BFS.scala 367:9]
  wire  _GEN_19 = _T & _T_16 ? io_in_bits_rdata[63:32] > 32'h0 : _GEN_18; // @[BFS.scala 370:72 BFS.scala 374:13]
  wire  keep_2 = _T & io_in_bits_rid[5] ? num_regfile_io_dataOut[63:32] > 32'h2 : _GEN_19; // @[BFS.scala 368:65 BFS.scala 369:11]
  wire  _GEN_21 = _T_8 & num > 32'h3; // @[BFS.scala 376:94 BFS.scala 377:11 BFS.scala 367:9]
  wire  _GEN_22 = _T & _T_16 ? io_in_bits_rdata[63:32] > 32'h1 : _GEN_21; // @[BFS.scala 370:72 BFS.scala 374:13]
  wire  keep_3 = _T & io_in_bits_rid[5] ? num_regfile_io_dataOut[63:32] > 32'h3 : _GEN_22; // @[BFS.scala 368:65 BFS.scala 369:11]
  wire [1:0] io_xbar_out_bits_tkeep_lo = {keep_1,keep_0}; // @[BFS.scala 384:40]
  wire [1:0] io_xbar_out_bits_tkeep_hi = {keep_3,keep_2}; // @[BFS.scala 384:40]
  wire [31:0] _edge_read_buffer_din_count_T_3 = io_in_bits_rdata[63:32] - 32'he; // @[BFS.scala 392:73]
  wire [31:0] _edge_read_buffer_din_index_T_4 = num_regfile_io_dataOut[31:0] + 32'h40; // @[BFS.scala 408:56]
  wire [31:0] _GEN_25 = num_regfile_io_dataOut[63:32] > 32'h40 ? _edge_read_buffer_din_index_T_4 : io_in_bits_rdata[31:0
    ]; // @[BFS.scala 404:85 BFS.scala 407:36 BFS.scala 393:30]
  wire [31:0] _GEN_30 = io_in_bits_rid[5] ? _GEN_25 : io_in_bits_rdata[31:0]; // @[BFS.scala 401:35 BFS.scala 393:30]
  wire [31:0] edge_read_buffer_din_index = _T_13 & _T ? _GEN_30 : io_in_bits_rdata[31:0]; // @[BFS.scala 399:64 BFS.scala 393:30]
  wire [4:0] _GEN_28 = io_in_bits_rid[5] ? io_in_bits_rid[4:0] : 5'h0; // @[BFS.scala 401:35 BFS.scala 403:36 BFS.scala 395:32]
  wire [4:0] _GEN_33 = _T_13 & _T ? _GEN_28 : 5'h0; // @[BFS.scala 399:64 BFS.scala 395:32]
  wire [5:0] edge_read_buffer_din_reg_ptr = {{1'd0}, _GEN_33}; // @[BFS.scala 389:34]
  wire [31:0] _edge_read_buffer_din_count_T_6 = num_regfile_io_dataOut[63:32] - 32'h40; // @[BFS.scala 406:50]
  wire [31:0] _GEN_24 = num_regfile_io_dataOut[63:32] > 32'h40 ? _edge_read_buffer_din_count_T_6 : 32'h0; // @[BFS.scala 404:85 BFS.scala 405:36 BFS.scala 410:36]
  wire [31:0] _GEN_26 = io_in_bits_rdata[63:32] < 32'he ? 32'h0 : _edge_read_buffer_din_count_T_3; // @[BFS.scala 413:66 BFS.scala 414:36 BFS.scala 392:30]
  wire [31:0] _GEN_29 = io_in_bits_rid[5] ? _GEN_24 : _GEN_26; // @[BFS.scala 401:35]
  wire [31:0] edge_read_buffer_din_count = _T_13 & _T ? _GEN_29 : _edge_read_buffer_din_count_T_3; // @[BFS.scala 399:64 BFS.scala 392:30]
  wire  _GEN_27 = io_in_bits_rid[5] ? 1'h0 : 1'h1; // @[BFS.scala 401:35 BFS.scala 402:35 BFS.scala 394:31]
  wire  edge_read_buffer_din_is_new = _T_13 & _T ? _GEN_27 : 1'h1; // @[BFS.scala 399:64 BFS.scala 394:31]
  wire [70:0] _edge_read_buffer_io_din_T = {edge_read_buffer_din_count,edge_read_buffer_din_is_new,
    edge_read_buffer_din_index,edge_read_buffer_din_reg_ptr}; // @[BFS.scala 398:57]
  wire [5:0] edge_read_buffer_dout_reg_ptr = edge_read_buffer__dout[5:0]; // @[BFS.scala 421:65]
  wire [31:0] edge_read_buffer_dout_index = edge_read_buffer__dout[37:6]; // @[BFS.scala 421:65]
  wire  edge_read_buffer_dout_is_new = edge_read_buffer__dout[38]; // @[BFS.scala 421:65]
  wire [31:0] edge_read_buffer_dout_count = edge_read_buffer__dout[70:39]; // @[BFS.scala 421:65]
  reg [3:0] cache_status; // @[BFS.scala 436:29]
  reg [5:0] init_seq; // @[BFS.scala 438:25]
  wire  _T_93 = cache_status == 4'h6; // @[BFS.scala 439:21]
  wire [5:0] _init_seq_T_1 = init_seq + 6'h1; // @[BFS.scala 440:26]
  reg [31:0] expand_index; // @[BFS.scala 442:29]
  reg [31:0] expand_count; // @[BFS.scala 443:29]
  reg [31:0] credit; // @[BFS.scala 444:23]
  wire  _T_100 = cache_status == 4'h0; // @[BFS.scala 449:27]
  wire  _T_103 = edge_read_buffer_dout_count == 32'h0; // @[BFS.scala 451:29]
  wire  _T_106 = edge_read_buffer_dout_count > 32'h40 & credit > 32'h4; // @[BFS.scala 454:65]
  wire [2:0] _GEN_37 = edge_read_buffer_dout_count > 32'h40 & credit > 32'h4 ? 3'h5 : 3'h2; // @[BFS.scala 454:99 BFS.scala 455:24 BFS.scala 459:24]
  wire [31:0] _GEN_38 = edge_read_buffer_dout_count > 32'h40 & credit > 32'h4 ? edge_read_buffer_dout_index :
    expand_index; // @[BFS.scala 454:99 BFS.scala 456:24 BFS.scala 442:29]
  wire [31:0] _GEN_39 = edge_read_buffer_dout_count > 32'h40 & credit > 32'h4 ? edge_read_buffer_dout_count :
    expand_count; // @[BFS.scala 454:99 BFS.scala 457:24 BFS.scala 443:29]
  wire [2:0] _GEN_40 = edge_read_buffer_dout_count == 32'h0 ? 3'h7 : _GEN_37; // @[BFS.scala 451:37 BFS.scala 452:22]
  wire [31:0] _GEN_41 = edge_read_buffer_dout_count == 32'h0 ? expand_index : _GEN_38; // @[BFS.scala 451:37 BFS.scala 442:29]
  wire [31:0] _GEN_42 = edge_read_buffer_dout_count == 32'h0 ? expand_count : _GEN_39; // @[BFS.scala 451:37 BFS.scala 443:29]
  wire [1:0] _GEN_43 = _T_106 ? 2'h1 : 2'h3; // @[BFS.scala 466:99 BFS.scala 467:24 BFS.scala 471:24]
  wire [2:0] _GEN_46 = _T_103 ? 3'h4 : {{1'd0}, _GEN_43}; // @[BFS.scala 463:37 BFS.scala 464:22]
  wire [2:0] _GEN_49 = edge_read_buffer_dout_is_new ? _GEN_40 : _GEN_46; // @[BFS.scala 450:50]
  wire [31:0] _GEN_50 = edge_read_buffer_dout_is_new ? _GEN_41 : _GEN_41; // @[BFS.scala 450:50]
  wire [31:0] _GEN_51 = edge_read_buffer_dout_is_new ? _GEN_42 : _GEN_42; // @[BFS.scala 450:50]
  wire  _T_111 = io_out_ready & io_out_valid; // @[BFS.scala 475:27]
  wire  _T_112 = cache_status == 4'h2; // @[BFS.scala 475:59]
  wire  _T_115 = cache_status == 4'h3; // @[BFS.scala 478:59]
  wire  _T_117 = cache_status == 4'h7; // @[BFS.scala 481:27]
  wire  _T_118 = cache_status == 4'h4; // @[BFS.scala 484:27]
  wire  _T_120 = cache_status == 4'h5; // @[BFS.scala 487:59]
  wire  _T_121 = _T_111 & cache_status == 4'h5; // @[BFS.scala 487:43]
  wire [31:0] _expand_index_T_1 = expand_index + 32'h40; // @[BFS.scala 488:34]
  wire [31:0] _expand_count_T_1 = expand_count - 32'h40; // @[BFS.scala 489:34]
  wire  _T_125 = credit <= 32'h4 | expand_count <= 32'h80; // @[BFS.scala 490:42]
  wire [3:0] _GEN_52 = credit <= 32'h4 | expand_count <= 32'h80 ? 4'h8 : cache_status; // @[BFS.scala 490:111 BFS.scala 491:20 BFS.scala 436:29]
  wire  _T_127 = cache_status == 4'h1; // @[BFS.scala 493:59]
  wire  _T_128 = _T_111 & cache_status == 4'h1; // @[BFS.scala 493:43]
  wire [3:0] _GEN_53 = _T_125 ? 4'h8 : 4'h5; // @[BFS.scala 496:111 BFS.scala 497:20 BFS.scala 499:20]
  wire  _T_134 = cache_status == 4'h8; // @[BFS.scala 501:59]
  wire  _T_135 = _T_111 & cache_status == 4'h8; // @[BFS.scala 501:43]
  wire [3:0] _GEN_54 = _T_111 & cache_status == 4'h8 ? 4'h0 : cache_status; // @[BFS.scala 501:83 BFS.scala 502:18 BFS.scala 436:29]
  wire [31:0] _GEN_56 = _T_111 & cache_status == 4'h1 ? _expand_index_T_1 : expand_index; // @[BFS.scala 493:91 BFS.scala 494:18 BFS.scala 442:29]
  wire [31:0] _GEN_57 = _T_111 & cache_status == 4'h1 ? _expand_count_T_1 : expand_count; // @[BFS.scala 493:91 BFS.scala 495:18 BFS.scala 443:29]
  wire [3:0] _GEN_58 = _T_111 & cache_status == 4'h1 ? _GEN_53 : _GEN_54; // @[BFS.scala 493:91]
  wire  _GEN_59 = _T_111 & cache_status == 4'h1 ? 1'h0 : _T_135; // @[BFS.scala 493:91 BFS.scala 397:29]
  wire [31:0] _GEN_60 = _T_111 & cache_status == 4'h5 ? _expand_index_T_1 : _GEN_56; // @[BFS.scala 487:91 BFS.scala 488:18]
  wire [31:0] _GEN_61 = _T_111 & cache_status == 4'h5 ? _expand_count_T_1 : _GEN_57; // @[BFS.scala 487:91 BFS.scala 489:18]
  wire [3:0] _GEN_62 = _T_111 & cache_status == 4'h5 ? _GEN_52 : _GEN_58; // @[BFS.scala 487:91]
  wire  _GEN_63 = _T_111 & cache_status == 4'h5 ? 1'h0 : _GEN_59; // @[BFS.scala 487:91 BFS.scala 397:29]
  wire [3:0] _GEN_64 = cache_status == 4'h4 ? 4'h0 : _GEN_62; // @[BFS.scala 484:51 BFS.scala 485:18]
  wire  _GEN_65 = cache_status == 4'h4 | _GEN_63; // @[BFS.scala 484:51 BFS.scala 486:31]
  wire [31:0] _GEN_66 = cache_status == 4'h4 ? expand_index : _GEN_60; // @[BFS.scala 484:51 BFS.scala 442:29]
  wire [31:0] _GEN_67 = cache_status == 4'h4 ? expand_count : _GEN_61; // @[BFS.scala 484:51 BFS.scala 443:29]
  wire [3:0] _GEN_68 = cache_status == 4'h7 ? 4'h0 : _GEN_64; // @[BFS.scala 481:55 BFS.scala 482:18]
  wire  _GEN_69 = cache_status == 4'h7 | _GEN_65; // @[BFS.scala 481:55 BFS.scala 483:31]
  wire [31:0] _GEN_70 = cache_status == 4'h7 ? expand_index : _GEN_66; // @[BFS.scala 481:55 BFS.scala 442:29]
  wire [31:0] _GEN_71 = cache_status == 4'h7 ? expand_count : _GEN_67; // @[BFS.scala 481:55 BFS.scala 443:29]
  wire [3:0] _GEN_72 = _T_111 & cache_status == 4'h3 ? 4'h0 : _GEN_68; // @[BFS.scala 478:87 BFS.scala 479:18]
  wire  _GEN_73 = _T_111 & cache_status == 4'h3 | _GEN_69; // @[BFS.scala 478:87 BFS.scala 480:31]
  wire [31:0] _GEN_74 = _T_111 & cache_status == 4'h3 ? expand_index : _GEN_70; // @[BFS.scala 478:87 BFS.scala 442:29]
  wire [31:0] _GEN_75 = _T_111 & cache_status == 4'h3 ? expand_count : _GEN_71; // @[BFS.scala 478:87 BFS.scala 443:29]
  wire [3:0] _GEN_76 = io_out_ready & io_out_valid & cache_status == 4'h2 ? 4'h0 : _GEN_72; // @[BFS.scala 475:84 BFS.scala 476:18]
  wire  _GEN_77 = io_out_ready & io_out_valid & cache_status == 4'h2 | _GEN_73; // @[BFS.scala 475:84 BFS.scala 477:31]
  wire [31:0] _GEN_78 = io_out_ready & io_out_valid & cache_status == 4'h2 ? expand_index : _GEN_74; // @[BFS.scala 475:84 BFS.scala 442:29]
  wire [31:0] _GEN_79 = io_out_ready & io_out_valid & cache_status == 4'h2 ? expand_count : _GEN_75; // @[BFS.scala 475:84 BFS.scala 443:29]
  wire  _GEN_83 = cache_status == 4'h0 & edge_read_buffer__valid ? 1'h0 : _GEN_77; // @[BFS.scala 449:77 BFS.scala 397:29]
  wire  _GEN_87 = _T_93 & init_seq == 6'h1f ? 1'h0 : _GEN_83; // @[BFS.scala 447:77 BFS.scala 397:29]
  wire  _num_vertex_T_2 = _T_134 & expand_count <= 32'h40; // @[BFS.scala 508:43]
  wire  _num_vertex_T_3 = edge_read_buffer_dout_count <= 32'h40; // @[BFS.scala 510:23]
  wire [31:0] _num_vertex_T_4 = _num_vertex_T_3 ? edge_read_buffer_dout_count : 32'h40; // @[Mux.scala 98:16]
  wire [31:0] num_vertex = _num_vertex_T_2 ? expand_count : _num_vertex_T_4; // @[Mux.scala 98:16]
  wire [31:0] _arlen_T_1 = {num_vertex[31:2], 2'h0}; // @[BFS.scala 512:63]
  wire [29:0] _arlen_T_6 = num_vertex[31:2] - 30'h1; // @[BFS.scala 514:57]
  wire [29:0] arlen = _arlen_T_1 < num_vertex ? num_vertex[31:2] : _arlen_T_6; // @[BFS.scala 512:18]
  wire [31:0] _io_out_bits_araddr_T_5 = _T_134 | _T_120 | _T_127 ? expand_index : edge_read_buffer_dout_index; // @[BFS.scala 517:11]
  wire [33:0] _GEN_131 = {_io_out_bits_araddr_T_5, 2'h0}; // @[BFS.scala 519:52]
  wire [34:0] _io_out_bits_araddr_T_6 = {{1'd0}, _GEN_131}; // @[BFS.scala 519:52]
  wire [63:0] _GEN_132 = {{29'd0}, _io_out_bits_araddr_T_6}; // @[BFS.scala 516:23]
  wire  _io_out_valid_T_4 = _T_112 | _T_115 | _T_134; // @[BFS.scala 520:100]
  wire  _io_out_bits_arsize_T = num_vertex <= 32'h1; // @[BFS.scala 527:23]
  wire  _io_out_bits_arsize_T_1 = num_vertex <= 32'h2; // @[BFS.scala 527:23]
  wire [2:0] _io_out_bits_arsize_T_2 = _io_out_bits_arsize_T_1 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  wire [4:0] io_out_bits_arid_lo = _T_112 | _T_120 | _T_134 ? free_queue_dout[4:0] : edge_read_buffer_dout_reg_ptr[4:0]; // @[BFS.scala 530:8]
  wire  _num_regfile_io_writeFlag_T_1 = free_queue_valid & io_out_ready & io_out_valid; // @[BFS.scala 547:71]
  wire [63:0] _num_regfile_io_dataIn_T = {edge_read_buffer_dout_count,edge_read_buffer_dout_index}; // @[Cat.scala 30:58]
  wire [38:0] _num_regfile_io_dataIn_T_2 = {7'h40,expand_index}; // @[Cat.scala 30:58]
  wire [63:0] _num_regfile_io_dataIn_T_4 = {expand_count,expand_index}; // @[Cat.scala 30:58]
  wire [5:0] _GEN_92 = _T_134 ? free_queue_dout : 6'h0; // @[BFS.scala 572:51 BFS.scala 573:25 BFS.scala 536:23]
  wire  _GEN_93 = _T_134 & _T_111; // @[BFS.scala 572:51 BFS.scala 574:25 BFS.scala 541:23]
  wire  _GEN_94 = _T_134 & _num_regfile_io_writeFlag_T_1; // @[BFS.scala 572:51 BFS.scala 575:30 BFS.scala 535:28]
  wire [63:0] _GEN_95 = _T_134 ? _num_regfile_io_dataIn_T_4 : 64'h0; // @[BFS.scala 572:51 BFS.scala 576:27 BFS.scala 537:25]
  wire [5:0] _GEN_96 = _T_127 ? edge_read_buffer_dout_reg_ptr : _GEN_92; // @[BFS.scala 567:59 BFS.scala 568:25]
  wire  _GEN_97 = _T_127 ? _T_111 : _GEN_94; // @[BFS.scala 567:59 BFS.scala 569:30]
  wire [63:0] _GEN_98 = _T_127 ? {{25'd0}, _num_regfile_io_dataIn_T_2} : _GEN_95; // @[BFS.scala 567:59 BFS.scala 570:27]
  wire  _GEN_99 = _T_127 ? 1'h0 : _GEN_93; // @[BFS.scala 567:59 BFS.scala 541:23]
  wire [5:0] _GEN_100 = _T_120 ? free_queue_dout : _GEN_96; // @[BFS.scala 561:59 BFS.scala 562:25]
  wire  _GEN_101 = _T_120 ? _T_111 : _GEN_99; // @[BFS.scala 561:59 BFS.scala 563:25]
  wire  _GEN_102 = _T_120 ? _num_regfile_io_writeFlag_T_1 : _GEN_97; // @[BFS.scala 561:59 BFS.scala 564:30]
  wire [63:0] _GEN_103 = _T_120 ? {{25'd0}, _num_regfile_io_dataIn_T_2} : _GEN_98; // @[BFS.scala 561:59 BFS.scala 565:27]
  wire [5:0] _GEN_104 = _T_93 ? init_seq : 6'h0; // @[BFS.scala 558:56 BFS.scala 559:23 BFS.scala 542:21]
  wire [5:0] _GEN_106 = _T_93 ? 6'h0 : _GEN_100; // @[BFS.scala 558:56 BFS.scala 536:23]
  wire  _GEN_107 = _T_93 ? 1'h0 : _GEN_101; // @[BFS.scala 558:56 BFS.scala 541:23]
  wire  _GEN_108 = _T_93 ? 1'h0 : _GEN_102; // @[BFS.scala 558:56 BFS.scala 535:28]
  wire [63:0] _GEN_109 = _T_93 ? 64'h0 : _GEN_103; // @[BFS.scala 558:56 BFS.scala 537:25]
  wire [5:0] _GEN_110 = _T_118 ? edge_read_buffer_dout_reg_ptr : _GEN_104; // @[BFS.scala 555:51 BFS.scala 556:23]
  wire  _GEN_111 = _T_118 | _T_93; // @[BFS.scala 555:51 BFS.scala 557:25]
  wire [5:0] _GEN_112 = _T_118 ? 6'h0 : _GEN_106; // @[BFS.scala 555:51 BFS.scala 536:23]
  wire  _GEN_113 = _T_118 ? 1'h0 : _GEN_107; // @[BFS.scala 555:51 BFS.scala 541:23]
  wire  _GEN_114 = _T_118 ? 1'h0 : _GEN_108; // @[BFS.scala 555:51 BFS.scala 535:28]
  wire [63:0] _GEN_115 = _T_118 ? 64'h0 : _GEN_109; // @[BFS.scala 555:51 BFS.scala 537:25]
  wire [5:0] _GEN_116 = _T_115 ? edge_read_buffer_dout_reg_ptr : _GEN_112; // @[BFS.scala 550:55 BFS.scala 551:25]
  wire  _GEN_117 = _T_115 ? _T_111 : _GEN_114; // @[BFS.scala 550:55 BFS.scala 552:30]
  wire [63:0] _GEN_118 = _T_115 ? _num_regfile_io_dataIn_T : _GEN_115; // @[BFS.scala 550:55 BFS.scala 553:27]
  wire [5:0] _GEN_119 = _T_115 ? 6'h0 : _GEN_110; // @[BFS.scala 550:55 BFS.scala 542:21]
  wire  _GEN_120 = _T_115 ? 1'h0 : _GEN_111; // @[BFS.scala 550:55 BFS.scala 543:23]
  wire  _GEN_121 = _T_115 ? 1'h0 : _GEN_113; // @[BFS.scala 550:55 BFS.scala 541:23]
  wire [5:0] _GEN_122 = _T_112 ? free_queue_dout : _GEN_116; // @[BFS.scala 544:46 BFS.scala 545:25]
  wire  _io_read_edge_fifo_empty_T = edge_read_buffer__data_count == 6'h0; // @[util.scala 211:19]
  wire  _credit_dec_T_6 = _T_121 | _T_128; // @[BFS.scala 582:97]
  wire  credit_dec = _credit_dec_T_6 | io_credit_dec; // @[BFS.scala 583:82]
  wire  _T_145 = cache_status != 4'h4; // @[BFS.scala 586:18]
  wire  _T_146 = credit_dec & cache_status != 4'h7 & _T_145; // @[BFS.scala 585:63]
  wire [31:0] _credit_T_1 = credit - 32'h1; // @[BFS.scala 587:22]
  wire  _T_151 = ~credit_dec & (_T_117 | _T_118); // @[BFS.scala 588:26]
  wire [31:0] _credit_T_3 = credit + 32'h1; // @[BFS.scala 590:22]
  regFile num_regfile ( // @[BFS.scala 341:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr)
  );
  meta_fifo edge_read_buffer_ ( // @[BFS.scala 387:32]
    .full(edge_read_buffer__full),
    .din(edge_read_buffer__din),
    .wr_en(edge_read_buffer__wr_en),
    .empty(edge_read_buffer__empty),
    .dout(edge_read_buffer__dout),
    .rd_en(edge_read_buffer__rd_en),
    .data_count(edge_read_buffer__data_count),
    .clk(edge_read_buffer__clk),
    .srst(edge_read_buffer__srst),
    .valid(edge_read_buffer__valid)
  );
  free_queue free_queue ( // @[BFS.scala 437:26]
    .full(free_queue_full),
    .din(free_queue_din),
    .wr_en(free_queue_wr_en),
    .empty(free_queue_empty),
    .dout(free_queue_dout),
    .rd_en(free_queue_rd_en),
    .data_count(free_queue_data_count),
    .clk(free_queue_clk),
    .srst(free_queue_srst),
    .valid(free_queue_valid)
  );
  assign io_in_ready = (~edge_read_buffer__full | status != 2'h0) & io_xbar_out_ready; // @[BFS.scala 418:84]
  assign io_out_valid = _io_out_valid_T_4 | _T_120 | _T_127; // @[BFS.scala 521:89]
  assign io_out_bits_araddr = io_edge_base_addr + _GEN_132; // @[BFS.scala 516:23]
  assign io_out_bits_arid = {1'h1,io_out_bits_arid_lo}; // @[Cat.scala 30:58]
  assign io_out_bits_arlen = arlen[7:0]; // @[BFS.scala 523:21]
  assign io_out_bits_arsize = _io_out_bits_arsize_T ? 3'h2 : _io_out_bits_arsize_T_2; // @[Mux.scala 98:16]
  assign io_xbar_out_valid = io_in_valid & io_in_ready; // @[BFS.scala 381:36]
  assign io_xbar_out_bits_tdata = io_in_bits_rdata; // @[BFS.scala 382:26]
  assign io_xbar_out_bits_tkeep = {io_xbar_out_bits_tkeep_hi,io_xbar_out_bits_tkeep_lo}; // @[BFS.scala 384:40]
  assign io_read_edge_fifo_empty = _io_read_edge_fifo_empty_T & _T_100; // @[BFS.scala 580:58]
  assign io_credit = credit[7:0]; // @[BFS.scala 592:13]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 338:21]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = _T_112 ? _num_regfile_io_dataIn_T : _GEN_118; // @[BFS.scala 544:46 BFS.scala 548:27]
  assign num_regfile_io_writeFlag = _T_112 ? free_queue_valid & io_out_ready & io_out_valid : _GEN_117; // @[BFS.scala 544:46 BFS.scala 547:30]
  assign num_regfile_io_rptr = io_in_bits_rid[4:0]; // @[BFS.scala 299:7]
  assign num_regfile_io_wptr = _GEN_122[4:0];
  assign edge_read_buffer__din = {{1'd0}, _edge_read_buffer_io_din_T}; // @[BFS.scala 398:57]
  assign edge_read_buffer__wr_en = _T_13 & _T; // @[BFS.scala 399:35]
  assign edge_read_buffer__rd_en = cache_status == 4'h9 & init_seq == 6'h0 ? 1'h0 : _GEN_87; // @[BFS.scala 445:60 BFS.scala 397:29]
  assign edge_read_buffer__clk = clock; // @[BFS.scala 390:42]
  assign edge_read_buffer__srst = reset; // @[BFS.scala 391:43]
  assign free_queue_din = _T_112 ? 6'h0 : _GEN_119; // @[BFS.scala 544:46 BFS.scala 542:21]
  assign free_queue_wr_en = _T_112 ? 1'h0 : _GEN_120; // @[BFS.scala 544:46 BFS.scala 543:23]
  assign free_queue_rd_en = _T_112 ? _T_111 : _GEN_121; // @[BFS.scala 544:46 BFS.scala 546:25]
  assign free_queue_clk = clock; // @[BFS.scala 539:36]
  assign free_queue_srst = reset; // @[BFS.scala 540:37]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 317:23]
      status <= 2'h0; // @[BFS.scala 317:23]
    end else if (status == 2'h0 & io_in_valid & io_in_ready) begin // @[BFS.scala 319:63]
      if (io_in_bits_rlast) begin // @[BFS.scala 320:36]
        status <= 2'h0; // @[BFS.scala 321:14]
      end else if (io_in_bits_rid[5]) begin // @[BFS.scala 322:41]
        status <= 2'h2; // @[BFS.scala 323:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 325:14]
      end
    end else if (_T_8 & io_in_valid & io_in_ready & io_in_bits_rlast) begin // @[BFS.scala 328:64]
      status <= 2'h0; // @[BFS.scala 329:12]
    end
    if (reset) begin // @[BFS.scala 318:20]
      num <= 32'h0; // @[BFS.scala 318:20]
    end else if (_T_2 & ~io_in_bits_rlast) begin // @[BFS.scala 343:65]
      if (io_in_bits_rid[5]) begin // @[BFS.scala 344:35]
        if (num_regfile_io_dataOut[63:32] > 32'h4) begin // @[BFS.scala 345:17]
          num <= _num_T_4;
        end else begin
          num <= 32'h0;
        end
      end else if (io_in_bits_rdata[63:32] > 32'h2) begin // @[BFS.scala 347:17]
        num <= _num_T_10;
      end else begin
        num <= 32'h0;
      end
    end else if (_T_6 & io_in_valid & io_in_ready) begin // @[BFS.scala 350:78]
      if (io_in_bits_rlast) begin // @[BFS.scala 351:36]
        num <= 32'h0; // @[BFS.scala 352:11]
      end else begin
        num <= _num_T_13; // @[BFS.scala 354:11]
      end
    end else if (_T_7 & io_in_valid & io_in_ready) begin // @[BFS.scala 356:83]
      num <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 331:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 331:35]
    end else if (io_signal) begin // @[BFS.scala 332:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 333:24]
    end else if (_T_17 & _T) begin // @[BFS.scala 335:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 336:24]
    end
    if (reset) begin // @[BFS.scala 436:29]
      cache_status <= 4'h9; // @[BFS.scala 436:29]
    end else if (cache_status == 4'h9 & init_seq == 6'h0) begin // @[BFS.scala 445:60]
      cache_status <= 4'h6; // @[BFS.scala 446:18]
    end else if (_T_93 & init_seq == 6'h1f) begin // @[BFS.scala 447:77]
      cache_status <= 4'h0; // @[BFS.scala 448:18]
    end else if (cache_status == 4'h0 & edge_read_buffer__valid) begin // @[BFS.scala 449:77]
      cache_status <= {{1'd0}, _GEN_49};
    end else begin
      cache_status <= _GEN_76;
    end
    if (reset) begin // @[BFS.scala 438:25]
      init_seq <= 6'h0; // @[BFS.scala 438:25]
    end else if (cache_status == 4'h6) begin // @[BFS.scala 439:50]
      init_seq <= _init_seq_T_1; // @[BFS.scala 440:14]
    end
    if (reset) begin // @[BFS.scala 442:29]
      expand_index <= 32'h0; // @[BFS.scala 442:29]
    end else if (!(cache_status == 4'h9 & init_seq == 6'h0)) begin // @[BFS.scala 445:60]
      if (!(_T_93 & init_seq == 6'h1f)) begin // @[BFS.scala 447:77]
        if (cache_status == 4'h0 & edge_read_buffer__valid) begin // @[BFS.scala 449:77]
          expand_index <= _GEN_50;
        end else begin
          expand_index <= _GEN_78;
        end
      end
    end
    if (reset) begin // @[BFS.scala 443:29]
      expand_count <= 32'h0; // @[BFS.scala 443:29]
    end else if (!(cache_status == 4'h9 & init_seq == 6'h0)) begin // @[BFS.scala 445:60]
      if (!(_T_93 & init_seq == 6'h1f)) begin // @[BFS.scala 447:77]
        if (cache_status == 4'h0 & edge_read_buffer__valid) begin // @[BFS.scala 449:77]
          expand_count <= _GEN_51;
        end else begin
          expand_count <= _GEN_79;
        end
      end
    end
    if (reset) begin // @[BFS.scala 444:23]
      credit <= 32'h20; // @[BFS.scala 444:23]
    end else if (_T_146) begin // @[BFS.scala 586:42]
      credit <= _credit_T_1; // @[BFS.scala 587:12]
    end else if (_T_151) begin // @[BFS.scala 589:43]
      credit <= _credit_T_3; // @[BFS.scala 590:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  status = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  num = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  cache_status = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  init_seq = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  expand_index = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  expand_count = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  credit = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AMBA_Arbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_araddr,
  input  [5:0]  io_in_0_bits_arid,
  input  [7:0]  io_in_0_bits_arlen,
  input  [2:0]  io_in_0_bits_arsize,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_araddr,
  input  [5:0]  io_in_1_bits_arid,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_araddr,
  output [5:0]  io_out_bits_arid,
  output [7:0]  io_out_bits_arlen,
  output [2:0]  io_out_bits_arsize
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  status; // @[util.scala 374:23]
  wire  grant_1 = ~io_in_0_valid; // @[util.scala 363:78]
  reg  grant_reg_0; // @[util.scala 376:26]
  reg  grant_reg_1; // @[util.scala 376:26]
  wire  _T = ~status; // @[util.scala 381:17]
  wire [2:0] _GEN_3 = io_in_0_valid ? io_in_0_bits_arsize : 3'h4; // @[util.scala 382:28 util.scala 384:21 util.scala 379:15]
  wire [7:0] _GEN_4 = io_in_0_valid ? io_in_0_bits_arlen : 8'h3; // @[util.scala 382:28 util.scala 384:21 util.scala 379:15]
  wire [5:0] _GEN_5 = io_in_0_valid ? io_in_0_bits_arid : io_in_1_bits_arid; // @[util.scala 382:28 util.scala 384:21 util.scala 379:15]
  wire [63:0] _GEN_6 = io_in_0_valid ? io_in_0_bits_araddr : io_in_1_bits_araddr; // @[util.scala 382:28 util.scala 384:21 util.scala 379:15]
  wire [2:0] _GEN_10 = grant_reg_0 ? io_in_0_bits_arsize : 3'h4; // @[util.scala 387:26 util.scala 389:21 util.scala 379:15]
  wire [7:0] _GEN_11 = grant_reg_0 ? io_in_0_bits_arlen : 8'h3; // @[util.scala 387:26 util.scala 389:21 util.scala 379:15]
  wire [5:0] _GEN_12 = grant_reg_0 ? io_in_0_bits_arid : io_in_1_bits_arid; // @[util.scala 387:26 util.scala 389:21 util.scala 379:15]
  wire [63:0] _GEN_13 = grant_reg_0 ? io_in_0_bits_araddr : io_in_1_bits_araddr; // @[util.scala 387:26 util.scala 389:21 util.scala 379:15]
  wire [2:0] _GEN_17 = status ? _GEN_10 : 3'h4; // @[util.scala 386:35 util.scala 379:15]
  wire [7:0] _GEN_18 = status ? _GEN_11 : 8'h3; // @[util.scala 386:35 util.scala 379:15]
  wire [5:0] _GEN_19 = status ? _GEN_12 : io_in_1_bits_arid; // @[util.scala 386:35 util.scala 379:15]
  wire [63:0] _GEN_20 = status ? _GEN_13 : io_in_1_bits_araddr; // @[util.scala 386:35 util.scala 379:15]
  wire  _T_8 = grant_1 & io_in_1_valid; // @[util.scala 396:24]
  wire  _GEN_28 = io_out_valid & io_out_ready & status ? 1'h0 : status; // @[util.scala 399:66 util.scala 400:12 util.scala 374:23]
  wire  _GEN_31 = (io_in_0_valid | io_in_1_valid) & _T & ~io_out_ready | _GEN_28; // @[util.scala 394:90 util.scala 398:12]
  assign io_in_0_ready = _T ? io_out_ready : grant_reg_0 & io_out_ready; // @[util.scala 403:20]
  assign io_in_1_ready = _T ? grant_1 & io_out_ready : grant_reg_1 & io_out_ready; // @[util.scala 403:20]
  assign io_out_valid = _T ? ~grant_1 | io_in_1_valid : ~grant_reg_1 | io_in_1_valid; // @[util.scala 405:22]
  assign io_out_bits_araddr = ~status ? _GEN_6 : _GEN_20; // @[util.scala 381:30]
  assign io_out_bits_arid = ~status ? _GEN_5 : _GEN_19; // @[util.scala 381:30]
  assign io_out_bits_arlen = ~status ? _GEN_4 : _GEN_18; // @[util.scala 381:30]
  assign io_out_bits_arsize = ~status ? _GEN_3 : _GEN_17; // @[util.scala 381:30]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 374:23]
      status <= 1'h0; // @[util.scala 374:23]
    end else begin
      status <= _GEN_31;
    end
    if (reset) begin // @[util.scala 376:26]
      grant_reg_0 <= 1'h0; // @[util.scala 376:26]
    end else if ((io_in_0_valid | io_in_1_valid) & _T & ~io_out_ready) begin // @[util.scala 394:90]
      grant_reg_0 <= io_in_0_valid; // @[util.scala 395:15]
    end
    if (reset) begin // @[util.scala 376:26]
      grant_reg_1 <= 1'h0; // @[util.scala 376:26]
    end else if ((io_in_0_valid | io_in_1_valid) & _T & ~io_out_ready) begin // @[util.scala 394:90]
      grant_reg_1 <= _T_8; // @[util.scala 395:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  status = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  grant_reg_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  grant_reg_1 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  output         io_xbar_out_bits_tlast,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  input          io_start,
  input  [31:0]  io_root,
  output         io_issue_sync,
  input  [4:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 633:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 633:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 633:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 633:34]
  wire  edge_cache_clock; // @[BFS.scala 640:26]
  wire  edge_cache_reset; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 640:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 640:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 640:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 640:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 640:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 640:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 640:26]
  wire  edge_cache_io_xbar_out_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_xbar_out_valid; // @[BFS.scala 640:26]
  wire [127:0] edge_cache_io_xbar_out_bits_tdata; // @[BFS.scala 640:26]
  wire [3:0] edge_cache_io_xbar_out_bits_tkeep; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 640:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 640:26]
  wire [7:0] edge_cache_io_credit; // @[BFS.scala 640:26]
  wire  edge_cache_io_credit_dec; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_traveled_edges; // @[BFS.scala 640:26]
  wire  edge_cache_io_signal; // @[BFS.scala 640:26]
  wire  arbi_clock; // @[BFS.scala 647:20]
  wire  arbi_reset; // @[BFS.scala 647:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 647:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 647:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 647:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 647:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 647:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 647:20]
  wire  arbi_io_out_ready; // @[BFS.scala 647:20]
  wire  arbi_io_out_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 647:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 647:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 647:20]
  wire  vertex_out_fifo_s_axis_aclk; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_aresetn; // @[BFS.scala 671:31]
  wire [127:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 671:31]
  wire [15:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 671:31]
  wire [127:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 671:31]
  wire [15:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 671:31]
  wire [31:0] vertex_out_fifo_axis_rd_data_count; // @[BFS.scala 671:31]
  reg [2:0] upward_status; // @[BFS.scala 629:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 630:30]
  reg [4:0] vertex_read_id; // @[BFS.scala 648:31]
  wire [4:0] _vertex_read_id_T_1 = vertex_read_id + 5'h1; // @[BFS.scala 650:38]
  wire [34:0] _arbi_io_in_1_bits_araddr_T_1 = {vertex_read_buffer_dout[30:2], 6'h0}; // @[BFS.scala 618:59]
  wire [63:0] _GEN_25 = {{29'd0}, _arbi_io_in_1_bits_araddr_T_1}; // @[BFS.scala 618:28]
  wire  _arbi_io_in_1_valid_T_3 = edge_cache_io_credit != 8'h0; // @[BFS.scala 655:26]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 661:104]
  wire [15:0] _io_xbar_out_bits_tkeep_T = vertex_out_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [127:0] _vertex_out_fifo_io_s_axis_tdata_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 128'h80000000 :
    edge_cache_io_xbar_out_bits_tdata; // @[Mux.scala 98:16]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 4'h1 :
    edge_cache_io_xbar_out_bits_tkeep; // @[Mux.scala 98:16]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_2 = io_start ? 4'h1 : _vertex_out_fifo_io_s_axis_tkeep_T_1; // @[Mux.scala 98:16]
  wire  _T_2 = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 689:81]
  reg [27:0] edge_fifo_ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_1 = edge_fifo_ready_counter + 28'h1; // @[Counter.scala 76:24]
  reg  syncRecv_0; // @[BFS.scala 693:25]
  reg  syncRecv_1; // @[BFS.scala 693:25]
  reg  syncRecv_2; // @[BFS.scala 693:25]
  reg  syncRecv_3; // @[BFS.scala 693:25]
  reg  syncRecv_4; // @[BFS.scala 693:25]
  wire  _GEN_4 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_6 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_8 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_10 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_12 = io_recv_sync[4] | syncRecv_4; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 703:34]
  wire [31:0] _T_11 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_15 = _T_11[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_25 = vertex_out_fifo_axis_rd_data_count == 32'h0; // @[util.scala 320:27]
  wire  _T_26 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_25; // @[BFS.scala 708:71]
  wire [2:0] _GEN_15 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 717:53 BFS.scala 718:19 BFS.scala 629:30]
  wire [2:0] _GEN_16 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3 & syncRecv_4) ? 3'h3 :
    _GEN_15; // @[BFS.scala 711:71]
  reg [27:0] ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_3 = ready_counter + 28'h1; // @[Counter.scala 76:24]
  wire  _T_38 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 724:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 728:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 730:36]
  wire  ar_ready_counter = 1'h0;
  vid_fifo vertex_read_buffer ( // @[BFS.scala 633:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 640:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_xbar_out_ready(edge_cache_io_xbar_out_ready),
    .io_xbar_out_valid(edge_cache_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(edge_cache_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(edge_cache_io_xbar_out_bits_tkeep),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_credit(edge_cache_io_credit),
    .io_credit_dec(edge_cache_io_credit_dec),
    .io_traveled_edges(edge_cache_io_traveled_edges),
    .io_signal(edge_cache_io_signal)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 647:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 671:31]
    .s_axis_aclk(vertex_out_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_out_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_out_fifo_axis_rd_data_count)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 652:13]
  assign io_ddr_r_ready = edge_cache_io_in_ready; // @[BFS.scala 643:20]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 638:52]
  assign io_xbar_out_valid = vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 675:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_xbar_out_bits_tlast = vertex_out_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_traveled_edges = edge_cache_io_traveled_edges; // @[BFS.scala 644:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 703:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 637:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 636:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 661:88]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 634:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 635:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = io_ddr_r_valid; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rdata = io_ddr_r_bits_rdata; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rid = io_ddr_r_bits_rid; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rlast = io_ddr_r_bits_rlast; // @[BFS.scala 643:20]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 662:17]
  assign edge_cache_io_xbar_out_ready = vertex_out_fifo_s_axis_tready; // @[BFS.scala 687:32]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 642:32]
  assign edge_cache_io_credit_dec = arbi_io_in_1_valid & arbi_io_in_1_ready; // @[BFS.scala 663:51]
  assign edge_cache_io_signal = io_signal; // @[BFS.scala 645:24]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 662:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & _arbi_io_in_1_valid_T_3; // @[BFS.scala 654:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_25; // @[BFS.scala 618:28]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 652:13]
  assign vertex_out_fifo_s_axis_aclk = clock; // @[BFS.scala 673:49]
  assign vertex_out_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 672:40]
  assign vertex_out_fifo_s_axis_tdata = io_start ? {{96'd0}, io_root} : _vertex_out_fifo_io_s_axis_tdata_T_1; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tvalid = edge_cache_io_xbar_out_valid | _vertex_read_buffer_io_rd_en_T_2 | io_start; // @[BFS.scala 677:109]
  assign vertex_out_fifo_s_axis_tkeep = {{12'd0}, _vertex_out_fifo_io_s_axis_tkeep_T_2}; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tlast = 1'h1; // @[BFS.scala 686:35]
  assign vertex_out_fifo_m_axis_tready = io_xbar_out_ready; // @[BFS.scala 676:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 629:30]
      upward_status <= 3'h0; // @[BFS.scala 629:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 704:57]
      upward_status <= 3'h1; // @[BFS.scala 705:19]
    end else if (upward_status == 3'h1 & (_T_15 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3 | syncRecv_4))
      ) begin // @[BFS.scala 706:105]
      upward_status <= 3'h2; // @[BFS.scala 707:19]
    end else if (_T_26 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 709:62]
      upward_status <= 3'h4; // @[BFS.scala 710:19]
    end else begin
      upward_status <= _GEN_16;
    end
    if (reset) begin // @[BFS.scala 630:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 630:30]
    end else if (!(_T_38 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 725:91]
      if (_T_38) begin // @[BFS.scala 727:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 728:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 729:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 730:19]
      end
    end
    if (reset) begin // @[BFS.scala 648:31]
      vertex_read_id <= 5'h0; // @[BFS.scala 648:31]
    end else if (arbi_io_in_1_valid & arbi_io_in_1_ready) begin // @[BFS.scala 649:51]
      vertex_read_id <= _vertex_read_id_T_1; // @[BFS.scala 650:20]
    end
    if (reset) begin // @[Counter.scala 60:40]
      edge_fifo_ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_2) begin // @[Counter.scala 118:17]
      edge_fifo_ready_counter <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_0 <= _GEN_4;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_1 <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_2 <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_3 <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_4 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_4 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_4 <= _GEN_12;
    end
    if (reset) begin // @[Counter.scala 60:40]
      ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_io_issue_sync_T) begin // @[Counter.scala 118:17]
      ready_counter <= _wrap_value_T_3; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  vertex_read_id = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  edge_fifo_ready_counter = _RAND_3[27:0];
  _RAND_4 = {1{`RANDOM}};
  syncRecv_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ready_counter = _RAND_9[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_1(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  output         io_xbar_out_bits_tlast,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [4:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 633:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 633:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 633:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 633:34]
  wire  edge_cache_clock; // @[BFS.scala 640:26]
  wire  edge_cache_reset; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 640:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 640:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 640:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 640:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 640:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 640:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 640:26]
  wire  edge_cache_io_xbar_out_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_xbar_out_valid; // @[BFS.scala 640:26]
  wire [127:0] edge_cache_io_xbar_out_bits_tdata; // @[BFS.scala 640:26]
  wire [3:0] edge_cache_io_xbar_out_bits_tkeep; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 640:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 640:26]
  wire [7:0] edge_cache_io_credit; // @[BFS.scala 640:26]
  wire  edge_cache_io_credit_dec; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_traveled_edges; // @[BFS.scala 640:26]
  wire  edge_cache_io_signal; // @[BFS.scala 640:26]
  wire  arbi_clock; // @[BFS.scala 647:20]
  wire  arbi_reset; // @[BFS.scala 647:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 647:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 647:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 647:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 647:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 647:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 647:20]
  wire  arbi_io_out_ready; // @[BFS.scala 647:20]
  wire  arbi_io_out_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 647:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 647:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 647:20]
  wire  vertex_out_fifo_s_axis_aclk; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_aresetn; // @[BFS.scala 671:31]
  wire [127:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 671:31]
  wire [15:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 671:31]
  wire [127:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 671:31]
  wire [15:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 671:31]
  wire [31:0] vertex_out_fifo_axis_rd_data_count; // @[BFS.scala 671:31]
  reg [2:0] upward_status; // @[BFS.scala 629:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 630:30]
  reg [4:0] vertex_read_id; // @[BFS.scala 648:31]
  wire [4:0] _vertex_read_id_T_1 = vertex_read_id + 5'h1; // @[BFS.scala 650:38]
  wire [34:0] _arbi_io_in_1_bits_araddr_T_1 = {vertex_read_buffer_dout[30:2], 6'h0}; // @[BFS.scala 618:59]
  wire [63:0] _GEN_25 = {{29'd0}, _arbi_io_in_1_bits_araddr_T_1}; // @[BFS.scala 618:28]
  wire  _arbi_io_in_1_valid_T_3 = edge_cache_io_credit != 8'h0; // @[BFS.scala 655:26]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 661:104]
  wire [15:0] _io_xbar_out_bits_tkeep_T = vertex_out_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 4'h1 :
    edge_cache_io_xbar_out_bits_tkeep; // @[Mux.scala 98:16]
  wire  _T_2 = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 689:81]
  reg [27:0] edge_fifo_ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_1 = edge_fifo_ready_counter + 28'h1; // @[Counter.scala 76:24]
  reg  syncRecv_0; // @[BFS.scala 693:25]
  reg  syncRecv_1; // @[BFS.scala 693:25]
  reg  syncRecv_2; // @[BFS.scala 693:25]
  reg  syncRecv_3; // @[BFS.scala 693:25]
  reg  syncRecv_4; // @[BFS.scala 693:25]
  wire  _GEN_4 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_6 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_8 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_10 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_12 = io_recv_sync[4] | syncRecv_4; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 703:34]
  wire [31:0] _T_11 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_15 = _T_11[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_25 = vertex_out_fifo_axis_rd_data_count == 32'h0; // @[util.scala 320:27]
  wire  _T_26 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_25; // @[BFS.scala 708:71]
  wire [2:0] _GEN_15 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 717:53 BFS.scala 718:19 BFS.scala 629:30]
  wire [2:0] _GEN_16 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3 & syncRecv_4) ? 3'h0 :
    _GEN_15; // @[BFS.scala 711:71]
  reg [27:0] ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_3 = ready_counter + 28'h1; // @[Counter.scala 76:24]
  wire  _T_38 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 724:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 728:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 730:36]
  wire  ar_ready_counter = 1'h0;
  vid_fifo vertex_read_buffer ( // @[BFS.scala 633:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 640:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_xbar_out_ready(edge_cache_io_xbar_out_ready),
    .io_xbar_out_valid(edge_cache_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(edge_cache_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(edge_cache_io_xbar_out_bits_tkeep),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_credit(edge_cache_io_credit),
    .io_credit_dec(edge_cache_io_credit_dec),
    .io_traveled_edges(edge_cache_io_traveled_edges),
    .io_signal(edge_cache_io_signal)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 647:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 671:31]
    .s_axis_aclk(vertex_out_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_out_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_out_fifo_axis_rd_data_count)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 652:13]
  assign io_ddr_r_ready = edge_cache_io_in_ready; // @[BFS.scala 643:20]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 638:52]
  assign io_xbar_out_valid = vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 675:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_xbar_out_bits_tlast = vertex_out_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_traveled_edges = edge_cache_io_traveled_edges; // @[BFS.scala 644:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 703:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 637:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 636:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 661:88]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 634:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 635:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = io_ddr_r_valid; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rdata = io_ddr_r_bits_rdata; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rid = io_ddr_r_bits_rid; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rlast = io_ddr_r_bits_rlast; // @[BFS.scala 643:20]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 662:17]
  assign edge_cache_io_xbar_out_ready = vertex_out_fifo_s_axis_tready; // @[BFS.scala 687:32]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 642:32]
  assign edge_cache_io_credit_dec = arbi_io_in_1_valid & arbi_io_in_1_ready; // @[BFS.scala 663:51]
  assign edge_cache_io_signal = io_signal; // @[BFS.scala 645:24]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 662:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & _arbi_io_in_1_valid_T_3; // @[BFS.scala 654:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_25; // @[BFS.scala 618:28]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 652:13]
  assign vertex_out_fifo_s_axis_aclk = clock; // @[BFS.scala 673:49]
  assign vertex_out_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 672:40]
  assign vertex_out_fifo_s_axis_tdata = _vertex_read_buffer_io_rd_en_T_2 ? 128'h80000000 :
    edge_cache_io_xbar_out_bits_tdata; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tvalid = edge_cache_io_xbar_out_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 677:68]
  assign vertex_out_fifo_s_axis_tkeep = {{12'd0}, _vertex_out_fifo_io_s_axis_tkeep_T_1}; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tlast = 1'h1; // @[BFS.scala 686:35]
  assign vertex_out_fifo_m_axis_tready = io_xbar_out_ready; // @[BFS.scala 676:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 629:30]
      upward_status <= 3'h0; // @[BFS.scala 629:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 704:57]
      upward_status <= 3'h1; // @[BFS.scala 705:19]
    end else if (upward_status == 3'h1 & (_T_15 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3 | syncRecv_4))
      ) begin // @[BFS.scala 706:105]
      upward_status <= 3'h2; // @[BFS.scala 707:19]
    end else if (_T_26 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 709:62]
      upward_status <= 3'h4; // @[BFS.scala 710:19]
    end else begin
      upward_status <= _GEN_16;
    end
    if (reset) begin // @[BFS.scala 630:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 630:30]
    end else if (!(_T_38 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 725:91]
      if (_T_38) begin // @[BFS.scala 727:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 728:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 729:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 730:19]
      end
    end
    if (reset) begin // @[BFS.scala 648:31]
      vertex_read_id <= 5'h0; // @[BFS.scala 648:31]
    end else if (arbi_io_in_1_valid & arbi_io_in_1_ready) begin // @[BFS.scala 649:51]
      vertex_read_id <= _vertex_read_id_T_1; // @[BFS.scala 650:20]
    end
    if (reset) begin // @[Counter.scala 60:40]
      edge_fifo_ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_2) begin // @[Counter.scala 118:17]
      edge_fifo_ready_counter <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_0 <= _GEN_4;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_1 <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_2 <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_3 <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_4 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_4 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_4 <= _GEN_12;
    end
    if (reset) begin // @[Counter.scala 60:40]
      ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_io_issue_sync_T) begin // @[Counter.scala 118:17]
      ready_counter <= _wrap_value_T_3; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  vertex_read_id = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  edge_fifo_ready_counter = _RAND_3[27:0];
  _RAND_4 = {1{`RANDOM}};
  syncRecv_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ready_counter = _RAND_9[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_2(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  output         io_xbar_out_bits_tlast,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [4:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 633:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 633:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 633:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 633:34]
  wire  edge_cache_clock; // @[BFS.scala 640:26]
  wire  edge_cache_reset; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 640:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 640:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 640:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 640:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 640:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 640:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 640:26]
  wire  edge_cache_io_xbar_out_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_xbar_out_valid; // @[BFS.scala 640:26]
  wire [127:0] edge_cache_io_xbar_out_bits_tdata; // @[BFS.scala 640:26]
  wire [3:0] edge_cache_io_xbar_out_bits_tkeep; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 640:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 640:26]
  wire [7:0] edge_cache_io_credit; // @[BFS.scala 640:26]
  wire  edge_cache_io_credit_dec; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_traveled_edges; // @[BFS.scala 640:26]
  wire  edge_cache_io_signal; // @[BFS.scala 640:26]
  wire  arbi_clock; // @[BFS.scala 647:20]
  wire  arbi_reset; // @[BFS.scala 647:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 647:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 647:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 647:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 647:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 647:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 647:20]
  wire  arbi_io_out_ready; // @[BFS.scala 647:20]
  wire  arbi_io_out_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 647:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 647:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 647:20]
  wire  vertex_out_fifo_s_axis_aclk; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_aresetn; // @[BFS.scala 671:31]
  wire [127:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 671:31]
  wire [15:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 671:31]
  wire [127:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 671:31]
  wire [15:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 671:31]
  wire [31:0] vertex_out_fifo_axis_rd_data_count; // @[BFS.scala 671:31]
  reg [2:0] upward_status; // @[BFS.scala 629:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 630:30]
  reg [4:0] vertex_read_id; // @[BFS.scala 648:31]
  wire [4:0] _vertex_read_id_T_1 = vertex_read_id + 5'h1; // @[BFS.scala 650:38]
  wire [34:0] _arbi_io_in_1_bits_araddr_T_1 = {vertex_read_buffer_dout[30:2], 6'h0}; // @[BFS.scala 618:59]
  wire [63:0] _GEN_25 = {{29'd0}, _arbi_io_in_1_bits_araddr_T_1}; // @[BFS.scala 618:28]
  wire  _arbi_io_in_1_valid_T_3 = edge_cache_io_credit != 8'h0; // @[BFS.scala 655:26]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 661:104]
  wire [15:0] _io_xbar_out_bits_tkeep_T = vertex_out_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 4'h1 :
    edge_cache_io_xbar_out_bits_tkeep; // @[Mux.scala 98:16]
  wire  _T_2 = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 689:81]
  reg [27:0] edge_fifo_ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_1 = edge_fifo_ready_counter + 28'h1; // @[Counter.scala 76:24]
  reg  syncRecv_0; // @[BFS.scala 693:25]
  reg  syncRecv_1; // @[BFS.scala 693:25]
  reg  syncRecv_2; // @[BFS.scala 693:25]
  reg  syncRecv_3; // @[BFS.scala 693:25]
  reg  syncRecv_4; // @[BFS.scala 693:25]
  wire  _GEN_4 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_6 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_8 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_10 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_12 = io_recv_sync[4] | syncRecv_4; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 703:34]
  wire [31:0] _T_11 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_15 = _T_11[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_25 = vertex_out_fifo_axis_rd_data_count == 32'h0; // @[util.scala 320:27]
  wire  _T_26 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_25; // @[BFS.scala 708:71]
  wire [2:0] _GEN_15 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 717:53 BFS.scala 718:19 BFS.scala 629:30]
  wire [2:0] _GEN_16 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3 & syncRecv_4) ? 3'h0 :
    _GEN_15; // @[BFS.scala 711:71]
  reg [27:0] ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_3 = ready_counter + 28'h1; // @[Counter.scala 76:24]
  wire  _T_38 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 724:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 728:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 730:36]
  wire  ar_ready_counter = 1'h0;
  vid_fifo vertex_read_buffer ( // @[BFS.scala 633:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 640:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_xbar_out_ready(edge_cache_io_xbar_out_ready),
    .io_xbar_out_valid(edge_cache_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(edge_cache_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(edge_cache_io_xbar_out_bits_tkeep),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_credit(edge_cache_io_credit),
    .io_credit_dec(edge_cache_io_credit_dec),
    .io_traveled_edges(edge_cache_io_traveled_edges),
    .io_signal(edge_cache_io_signal)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 647:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 671:31]
    .s_axis_aclk(vertex_out_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_out_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_out_fifo_axis_rd_data_count)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 652:13]
  assign io_ddr_r_ready = edge_cache_io_in_ready; // @[BFS.scala 643:20]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 638:52]
  assign io_xbar_out_valid = vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 675:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_xbar_out_bits_tlast = vertex_out_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_traveled_edges = edge_cache_io_traveled_edges; // @[BFS.scala 644:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 703:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 637:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 636:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 661:88]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 634:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 635:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = io_ddr_r_valid; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rdata = io_ddr_r_bits_rdata; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rid = io_ddr_r_bits_rid; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rlast = io_ddr_r_bits_rlast; // @[BFS.scala 643:20]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 662:17]
  assign edge_cache_io_xbar_out_ready = vertex_out_fifo_s_axis_tready; // @[BFS.scala 687:32]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 642:32]
  assign edge_cache_io_credit_dec = arbi_io_in_1_valid & arbi_io_in_1_ready; // @[BFS.scala 663:51]
  assign edge_cache_io_signal = io_signal; // @[BFS.scala 645:24]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 662:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & _arbi_io_in_1_valid_T_3; // @[BFS.scala 654:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_25; // @[BFS.scala 618:28]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 652:13]
  assign vertex_out_fifo_s_axis_aclk = clock; // @[BFS.scala 673:49]
  assign vertex_out_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 672:40]
  assign vertex_out_fifo_s_axis_tdata = _vertex_read_buffer_io_rd_en_T_2 ? 128'h80000000 :
    edge_cache_io_xbar_out_bits_tdata; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tvalid = edge_cache_io_xbar_out_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 677:68]
  assign vertex_out_fifo_s_axis_tkeep = {{12'd0}, _vertex_out_fifo_io_s_axis_tkeep_T_1}; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tlast = 1'h1; // @[BFS.scala 686:35]
  assign vertex_out_fifo_m_axis_tready = io_xbar_out_ready; // @[BFS.scala 676:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 629:30]
      upward_status <= 3'h0; // @[BFS.scala 629:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 704:57]
      upward_status <= 3'h1; // @[BFS.scala 705:19]
    end else if (upward_status == 3'h1 & (_T_15 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3 | syncRecv_4))
      ) begin // @[BFS.scala 706:105]
      upward_status <= 3'h2; // @[BFS.scala 707:19]
    end else if (_T_26 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 709:62]
      upward_status <= 3'h4; // @[BFS.scala 710:19]
    end else begin
      upward_status <= _GEN_16;
    end
    if (reset) begin // @[BFS.scala 630:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 630:30]
    end else if (!(_T_38 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 725:91]
      if (_T_38) begin // @[BFS.scala 727:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 728:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 729:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 730:19]
      end
    end
    if (reset) begin // @[BFS.scala 648:31]
      vertex_read_id <= 5'h0; // @[BFS.scala 648:31]
    end else if (arbi_io_in_1_valid & arbi_io_in_1_ready) begin // @[BFS.scala 649:51]
      vertex_read_id <= _vertex_read_id_T_1; // @[BFS.scala 650:20]
    end
    if (reset) begin // @[Counter.scala 60:40]
      edge_fifo_ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_2) begin // @[Counter.scala 118:17]
      edge_fifo_ready_counter <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_0 <= _GEN_4;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_1 <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_2 <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_3 <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_4 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_4 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_4 <= _GEN_12;
    end
    if (reset) begin // @[Counter.scala 60:40]
      ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_io_issue_sync_T) begin // @[Counter.scala 118:17]
      ready_counter <= _wrap_value_T_3; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  vertex_read_id = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  edge_fifo_ready_counter = _RAND_3[27:0];
  _RAND_4 = {1{`RANDOM}};
  syncRecv_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ready_counter = _RAND_9[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_3(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  output         io_xbar_out_bits_tlast,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [4:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 633:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 633:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 633:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 633:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 633:34]
  wire  edge_cache_clock; // @[BFS.scala 640:26]
  wire  edge_cache_reset; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 640:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 640:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 640:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 640:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 640:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 640:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 640:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 640:26]
  wire  edge_cache_io_xbar_out_ready; // @[BFS.scala 640:26]
  wire  edge_cache_io_xbar_out_valid; // @[BFS.scala 640:26]
  wire [127:0] edge_cache_io_xbar_out_bits_tdata; // @[BFS.scala 640:26]
  wire [3:0] edge_cache_io_xbar_out_bits_tkeep; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 640:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 640:26]
  wire [7:0] edge_cache_io_credit; // @[BFS.scala 640:26]
  wire  edge_cache_io_credit_dec; // @[BFS.scala 640:26]
  wire [63:0] edge_cache_io_traveled_edges; // @[BFS.scala 640:26]
  wire  edge_cache_io_signal; // @[BFS.scala 640:26]
  wire  arbi_clock; // @[BFS.scala 647:20]
  wire  arbi_reset; // @[BFS.scala 647:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 647:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 647:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 647:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 647:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 647:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 647:20]
  wire  arbi_io_out_ready; // @[BFS.scala 647:20]
  wire  arbi_io_out_valid; // @[BFS.scala 647:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 647:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 647:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 647:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 647:20]
  wire  vertex_out_fifo_s_axis_aclk; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_aresetn; // @[BFS.scala 671:31]
  wire [127:0] vertex_out_fifo_s_axis_tdata; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tvalid; // @[BFS.scala 671:31]
  wire [15:0] vertex_out_fifo_s_axis_tkeep; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tready; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_s_axis_tlast; // @[BFS.scala 671:31]
  wire [127:0] vertex_out_fifo_m_axis_tdata; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 671:31]
  wire [15:0] vertex_out_fifo_m_axis_tkeep; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tready; // @[BFS.scala 671:31]
  wire  vertex_out_fifo_m_axis_tlast; // @[BFS.scala 671:31]
  wire [31:0] vertex_out_fifo_axis_rd_data_count; // @[BFS.scala 671:31]
  reg [2:0] upward_status; // @[BFS.scala 629:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 630:30]
  reg [4:0] vertex_read_id; // @[BFS.scala 648:31]
  wire [4:0] _vertex_read_id_T_1 = vertex_read_id + 5'h1; // @[BFS.scala 650:38]
  wire [34:0] _arbi_io_in_1_bits_araddr_T_1 = {vertex_read_buffer_dout[30:2], 6'h0}; // @[BFS.scala 618:59]
  wire [63:0] _GEN_25 = {{29'd0}, _arbi_io_in_1_bits_araddr_T_1}; // @[BFS.scala 618:28]
  wire  _arbi_io_in_1_valid_T_3 = edge_cache_io_credit != 8'h0; // @[BFS.scala 655:26]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 661:104]
  wire [15:0] _io_xbar_out_bits_tkeep_T = vertex_out_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [3:0] _vertex_out_fifo_io_s_axis_tkeep_T_1 = _vertex_read_buffer_io_rd_en_T_2 ? 4'h1 :
    edge_cache_io_xbar_out_bits_tkeep; // @[Mux.scala 98:16]
  wire  _T_2 = ~vertex_out_fifo_s_axis_tready; // @[BFS.scala 689:81]
  reg [27:0] edge_fifo_ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_1 = edge_fifo_ready_counter + 28'h1; // @[Counter.scala 76:24]
  reg  syncRecv_0; // @[BFS.scala 693:25]
  reg  syncRecv_1; // @[BFS.scala 693:25]
  reg  syncRecv_2; // @[BFS.scala 693:25]
  reg  syncRecv_3; // @[BFS.scala 693:25]
  reg  syncRecv_4; // @[BFS.scala 693:25]
  wire  _GEN_4 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_6 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_8 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_10 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _GEN_12 = io_recv_sync[4] | syncRecv_4; // @[BFS.scala 698:34 BFS.scala 699:11 BFS.scala 693:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 703:34]
  wire [31:0] _T_11 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_15 = _T_11[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_25 = vertex_out_fifo_axis_rd_data_count == 32'h0; // @[util.scala 320:27]
  wire  _T_26 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_25; // @[BFS.scala 708:71]
  wire [2:0] _GEN_15 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 717:53 BFS.scala 718:19 BFS.scala 629:30]
  wire [2:0] _GEN_16 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3 & syncRecv_4) ? 3'h0 :
    _GEN_15; // @[BFS.scala 711:71]
  reg [27:0] ready_counter; // @[Counter.scala 60:40]
  wire [27:0] _wrap_value_T_3 = ready_counter + 28'h1; // @[Counter.scala 76:24]
  wire  _T_38 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 724:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 728:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 730:36]
  wire  ar_ready_counter = 1'h0;
  vid_fifo vertex_read_buffer ( // @[BFS.scala 633:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 640:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_xbar_out_ready(edge_cache_io_xbar_out_ready),
    .io_xbar_out_valid(edge_cache_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(edge_cache_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(edge_cache_io_xbar_out_bits_tkeep),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_credit(edge_cache_io_credit),
    .io_credit_dec(edge_cache_io_credit_dec),
    .io_traveled_edges(edge_cache_io_traveled_edges),
    .io_signal(edge_cache_io_signal)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 647:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 671:31]
    .s_axis_aclk(vertex_out_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_out_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_out_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_out_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_out_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_out_fifo_s_axis_tready),
    .s_axis_tlast(vertex_out_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_out_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_out_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_out_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_out_fifo_m_axis_tready),
    .m_axis_tlast(vertex_out_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_out_fifo_axis_rd_data_count)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 652:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 652:13]
  assign io_ddr_r_ready = edge_cache_io_in_ready; // @[BFS.scala 643:20]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 638:52]
  assign io_xbar_out_valid = vertex_out_fifo_m_axis_tvalid; // @[BFS.scala 675:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_xbar_out_bits_tlast = vertex_out_fifo_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_traveled_edges = edge_cache_io_traveled_edges; // @[BFS.scala 644:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 703:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 637:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 636:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 661:88]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 634:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 635:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = io_ddr_r_valid; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rdata = io_ddr_r_bits_rdata; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rid = io_ddr_r_bits_rid; // @[BFS.scala 643:20]
  assign edge_cache_io_in_bits_rlast = io_ddr_r_bits_rlast; // @[BFS.scala 643:20]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 662:17]
  assign edge_cache_io_xbar_out_ready = vertex_out_fifo_s_axis_tready; // @[BFS.scala 687:32]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 642:32]
  assign edge_cache_io_credit_dec = arbi_io_in_1_valid & arbi_io_in_1_ready; // @[BFS.scala 663:51]
  assign edge_cache_io_signal = io_signal; // @[BFS.scala 645:24]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 662:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 662:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & _arbi_io_in_1_valid_T_3; // @[BFS.scala 654:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_25; // @[BFS.scala 618:28]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 652:13]
  assign vertex_out_fifo_s_axis_aclk = clock; // @[BFS.scala 673:49]
  assign vertex_out_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 672:40]
  assign vertex_out_fifo_s_axis_tdata = _vertex_read_buffer_io_rd_en_T_2 ? 128'h80000000 :
    edge_cache_io_xbar_out_bits_tdata; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tvalid = edge_cache_io_xbar_out_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 677:68]
  assign vertex_out_fifo_s_axis_tkeep = {{12'd0}, _vertex_out_fifo_io_s_axis_tkeep_T_1}; // @[Mux.scala 98:16]
  assign vertex_out_fifo_s_axis_tlast = 1'h1; // @[BFS.scala 686:35]
  assign vertex_out_fifo_m_axis_tready = io_xbar_out_ready; // @[BFS.scala 676:36]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 629:30]
      upward_status <= 3'h0; // @[BFS.scala 629:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 704:57]
      upward_status <= 3'h1; // @[BFS.scala 705:19]
    end else if (upward_status == 3'h1 & (_T_15 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3 | syncRecv_4))
      ) begin // @[BFS.scala 706:105]
      upward_status <= 3'h2; // @[BFS.scala 707:19]
    end else if (_T_26 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 709:62]
      upward_status <= 3'h4; // @[BFS.scala 710:19]
    end else begin
      upward_status <= _GEN_16;
    end
    if (reset) begin // @[BFS.scala 630:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 630:30]
    end else if (!(_T_38 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 725:91]
      if (_T_38) begin // @[BFS.scala 727:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 728:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 729:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 730:19]
      end
    end
    if (reset) begin // @[BFS.scala 648:31]
      vertex_read_id <= 5'h0; // @[BFS.scala 648:31]
    end else if (arbi_io_in_1_valid & arbi_io_in_1_ready) begin // @[BFS.scala 649:51]
      vertex_read_id <= _vertex_read_id_T_1; // @[BFS.scala 650:20]
    end
    if (reset) begin // @[Counter.scala 60:40]
      edge_fifo_ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_T_2) begin // @[Counter.scala 118:17]
      edge_fifo_ready_counter <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_0 <= _GEN_4;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_1 <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_2 <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_3 <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 693:25]
      syncRecv_4 <= 1'h0; // @[BFS.scala 693:25]
    end else if (io_signal) begin // @[BFS.scala 696:22]
      syncRecv_4 <= 1'h0; // @[BFS.scala 697:11]
    end else begin
      syncRecv_4 <= _GEN_12;
    end
    if (reset) begin // @[Counter.scala 60:40]
      ready_counter <= 28'h0; // @[Counter.scala 60:40]
    end else if (_io_issue_sync_T) begin // @[Counter.scala 118:17]
      ready_counter <= _wrap_value_T_3; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  vertex_read_id = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  edge_fifo_ready_counter = _RAND_3[27:0];
  _RAND_4 = {1{`RANDOM}};
  syncRecv_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ready_counter = _RAND_9[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_data_collector(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [511:0] io_in_bits_tdata,
  input  [15:0]  io_in_bits_tkeep,
  input          io_out_ready,
  output         io_out_valid,
  output [511:0] io_out_bits_tdata,
  output [15:0]  io_out_bits_tkeep,
  output         io_out_bits_tlast,
  input          io_flush,
  output         io_empty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  in_aclk; // @[bfs_remote.scala 19:18]
  wire  in_aresetn; // @[bfs_remote.scala 19:18]
  wire [511:0] in_s_axis_tdata; // @[bfs_remote.scala 19:18]
  wire  in_s_axis_tvalid; // @[bfs_remote.scala 19:18]
  wire [63:0] in_s_axis_tkeep; // @[bfs_remote.scala 19:18]
  wire  in_s_axis_tready; // @[bfs_remote.scala 19:18]
  wire  in_s_axis_tlast; // @[bfs_remote.scala 19:18]
  wire [511:0] in_m_axis_tdata; // @[bfs_remote.scala 19:18]
  wire  in_m_axis_tvalid; // @[bfs_remote.scala 19:18]
  wire [63:0] in_m_axis_tkeep; // @[bfs_remote.scala 19:18]
  wire  in_m_axis_tready; // @[bfs_remote.scala 19:18]
  wire  in_m_axis_tlast; // @[bfs_remote.scala 19:18]
  wire  sorted_in_aclk; // @[bfs_remote.scala 43:25]
  wire  sorted_in_aresetn; // @[bfs_remote.scala 43:25]
  wire [511:0] sorted_in_s_axis_tdata; // @[bfs_remote.scala 43:25]
  wire  sorted_in_s_axis_tvalid; // @[bfs_remote.scala 43:25]
  wire [63:0] sorted_in_s_axis_tkeep; // @[bfs_remote.scala 43:25]
  wire  sorted_in_s_axis_tready; // @[bfs_remote.scala 43:25]
  wire  sorted_in_s_axis_tlast; // @[bfs_remote.scala 43:25]
  wire [511:0] sorted_in_m_axis_tdata; // @[bfs_remote.scala 43:25]
  wire  sorted_in_m_axis_tvalid; // @[bfs_remote.scala 43:25]
  wire [63:0] sorted_in_m_axis_tkeep; // @[bfs_remote.scala 43:25]
  wire  sorted_in_m_axis_tready; // @[bfs_remote.scala 43:25]
  wire  sorted_in_m_axis_tlast; // @[bfs_remote.scala 43:25]
  wire  mid_aclk; // @[bfs_remote.scala 55:19]
  wire  mid_aresetn; // @[bfs_remote.scala 55:19]
  wire [1023:0] mid_s_axis_tdata; // @[bfs_remote.scala 55:19]
  wire  mid_s_axis_tvalid; // @[bfs_remote.scala 55:19]
  wire [127:0] mid_s_axis_tkeep; // @[bfs_remote.scala 55:19]
  wire  mid_s_axis_tready; // @[bfs_remote.scala 55:19]
  wire  mid_s_axis_tlast; // @[bfs_remote.scala 55:19]
  wire [1023:0] mid_m_axis_tdata; // @[bfs_remote.scala 55:19]
  wire  mid_m_axis_tvalid; // @[bfs_remote.scala 55:19]
  wire [127:0] mid_m_axis_tkeep; // @[bfs_remote.scala 55:19]
  wire  mid_m_axis_tready; // @[bfs_remote.scala 55:19]
  wire  mid_m_axis_tlast; // @[bfs_remote.scala 55:19]
  wire  out_aclk; // @[bfs_remote.scala 86:19]
  wire  out_aresetn; // @[bfs_remote.scala 86:19]
  wire [511:0] out_s_axis_tdata; // @[bfs_remote.scala 86:19]
  wire  out_s_axis_tvalid; // @[bfs_remote.scala 86:19]
  wire [63:0] out_s_axis_tkeep; // @[bfs_remote.scala 86:19]
  wire  out_s_axis_tready; // @[bfs_remote.scala 86:19]
  wire  out_s_axis_tlast; // @[bfs_remote.scala 86:19]
  wire [511:0] out_m_axis_tdata; // @[bfs_remote.scala 86:19]
  wire  out_m_axis_tvalid; // @[bfs_remote.scala 86:19]
  wire [63:0] out_m_axis_tkeep; // @[bfs_remote.scala 86:19]
  wire  out_m_axis_tready; // @[bfs_remote.scala 86:19]
  wire  out_m_axis_tlast; // @[bfs_remote.scala 86:19]
  wire  _in_count_T_18 = in_m_axis_tkeep[0] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire  _in_count_T_56 = in_m_axis_tkeep[1] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE = {{7'd0}, _in_count_T_18}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] _in_count_WIRE_1 = {{7'd0}, _in_count_T_56}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_1 = _in_count_WIRE + _in_count_WIRE_1; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_114 = in_m_axis_tkeep[2] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_4 = {{7'd0}, _in_count_T_114}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_2 = in_count_1 + _in_count_WIRE_4; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_193 = in_m_axis_tkeep[3] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_8 = {{7'd0}, _in_count_T_193}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_3 = in_count_2 + _in_count_WIRE_8; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_293 = in_m_axis_tkeep[4] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_13 = {{7'd0}, _in_count_T_293}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_4 = in_count_3 + _in_count_WIRE_13; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_414 = in_m_axis_tkeep[5] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_19 = {{7'd0}, _in_count_T_414}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_5 = in_count_4 + _in_count_WIRE_19; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_556 = in_m_axis_tkeep[6] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_26 = {{7'd0}, _in_count_T_556}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_6 = in_count_5 + _in_count_WIRE_26; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_719 = in_m_axis_tkeep[7] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_34 = {{7'd0}, _in_count_T_719}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_7 = in_count_6 + _in_count_WIRE_34; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_903 = in_m_axis_tkeep[8] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_43 = {{7'd0}, _in_count_T_903}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_8 = in_count_7 + _in_count_WIRE_43; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_1108 = in_m_axis_tkeep[9] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_53 = {{7'd0}, _in_count_T_1108}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_9 = in_count_8 + _in_count_WIRE_53; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_1334 = in_m_axis_tkeep[10] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_64 = {{7'd0}, _in_count_T_1334}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_10 = in_count_9 + _in_count_WIRE_64; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_1581 = in_m_axis_tkeep[11] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_76 = {{7'd0}, _in_count_T_1581}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_11 = in_count_10 + _in_count_WIRE_76; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_1849 = in_m_axis_tkeep[12] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_89 = {{7'd0}, _in_count_T_1849}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_12 = in_count_11 + _in_count_WIRE_89; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_2138 = in_m_axis_tkeep[13] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_103 = {{7'd0}, _in_count_T_2138}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_13 = in_count_12 + _in_count_WIRE_103; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_2448 = in_m_axis_tkeep[14] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_118 = {{7'd0}, _in_count_T_2448}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_14 = in_count_13 + _in_count_WIRE_118; // @[bfs_remote.scala 28:151]
  wire  _in_count_T_2779 = in_m_axis_tkeep[15] & in_m_axis_tvalid; // @[bfs_remote.scala 28:89]
  wire [7:0] _in_count_WIRE_134 = {{7'd0}, _in_count_T_2779}; // @[bfs_remote.scala 28:130 bfs_remote.scala 28:130]
  wire [7:0] in_count_15 = in_count_14 + _in_count_WIRE_134; // @[bfs_remote.scala 28:151]
  wire  _in_data_0_tdata_T_2 = 8'h1 == _in_count_WIRE; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_6 = 8'h1 == in_count_1; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_10 = 8'h1 == in_count_2; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_14 = 8'h1 == in_count_3; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_18 = 8'h1 == in_count_4; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_22 = 8'h1 == in_count_5; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_26 = 8'h1 == in_count_6; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_30 = 8'h1 == in_count_7; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_34 = 8'h1 == in_count_8; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_38 = 8'h1 == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_42 = 8'h1 == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_46 = 8'h1 == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_50 = 8'h1 == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_54 = 8'h1 == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_58 = 8'h1 == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_0_tdata_T_62 = 8'h1 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_0_tdata_T_64 = _in_data_0_tdata_T_62 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_65 = _in_data_0_tdata_T_58 ? in_m_axis_tdata[479:448] : _in_data_0_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_66 = _in_data_0_tdata_T_54 ? in_m_axis_tdata[447:416] : _in_data_0_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_67 = _in_data_0_tdata_T_50 ? in_m_axis_tdata[415:384] : _in_data_0_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_68 = _in_data_0_tdata_T_46 ? in_m_axis_tdata[383:352] : _in_data_0_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_69 = _in_data_0_tdata_T_42 ? in_m_axis_tdata[351:320] : _in_data_0_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_70 = _in_data_0_tdata_T_38 ? in_m_axis_tdata[319:288] : _in_data_0_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_71 = _in_data_0_tdata_T_34 ? in_m_axis_tdata[287:256] : _in_data_0_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_72 = _in_data_0_tdata_T_30 ? in_m_axis_tdata[255:224] : _in_data_0_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_73 = _in_data_0_tdata_T_26 ? in_m_axis_tdata[223:192] : _in_data_0_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_74 = _in_data_0_tdata_T_22 ? in_m_axis_tdata[191:160] : _in_data_0_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_75 = _in_data_0_tdata_T_18 ? in_m_axis_tdata[159:128] : _in_data_0_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_76 = _in_data_0_tdata_T_14 ? in_m_axis_tdata[127:96] : _in_data_0_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_77 = _in_data_0_tdata_T_10 ? in_m_axis_tdata[95:64] : _in_data_0_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _in_data_0_tdata_T_78 = _in_data_0_tdata_T_6 ? in_m_axis_tdata[63:32] : _in_data_0_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] in_data_0_tdata = _in_data_0_tdata_T_2 ? in_m_axis_tdata[31:0] : _in_data_0_tdata_T_78; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_65 = _in_data_0_tdata_T_58 ? in_m_axis_tkeep[14] : _in_data_0_tdata_T_62 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_66 = _in_data_0_tdata_T_54 ? in_m_axis_tkeep[13] : _in_data_0_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_67 = _in_data_0_tdata_T_50 ? in_m_axis_tkeep[12] : _in_data_0_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_68 = _in_data_0_tdata_T_46 ? in_m_axis_tkeep[11] : _in_data_0_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_69 = _in_data_0_tdata_T_42 ? in_m_axis_tkeep[10] : _in_data_0_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_70 = _in_data_0_tdata_T_38 ? in_m_axis_tkeep[9] : _in_data_0_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_71 = _in_data_0_tdata_T_34 ? in_m_axis_tkeep[8] : _in_data_0_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_72 = _in_data_0_tdata_T_30 ? in_m_axis_tkeep[7] : _in_data_0_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_73 = _in_data_0_tdata_T_26 ? in_m_axis_tkeep[6] : _in_data_0_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_74 = _in_data_0_tdata_T_22 ? in_m_axis_tkeep[5] : _in_data_0_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_75 = _in_data_0_tdata_T_18 ? in_m_axis_tkeep[4] : _in_data_0_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_76 = _in_data_0_tdata_T_14 ? in_m_axis_tkeep[3] : _in_data_0_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_77 = _in_data_0_tdata_T_10 ? in_m_axis_tkeep[2] : _in_data_0_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _in_data_0_tkeep_T_78 = _in_data_0_tdata_T_6 ? in_m_axis_tkeep[1] : _in_data_0_tkeep_T_77; // @[Mux.scala 98:16]
  wire  in_data_0_tkeep = _in_data_0_tdata_T_2 ? in_m_axis_tkeep[0] : _in_data_0_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _in_data_1_tdata_T_2 = 8'h2 == in_count_1; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_6 = 8'h2 == in_count_2; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_10 = 8'h2 == in_count_3; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_14 = 8'h2 == in_count_4; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_18 = 8'h2 == in_count_5; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_22 = 8'h2 == in_count_6; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_26 = 8'h2 == in_count_7; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_30 = 8'h2 == in_count_8; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_34 = 8'h2 == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_38 = 8'h2 == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_42 = 8'h2 == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_46 = 8'h2 == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_50 = 8'h2 == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_54 = 8'h2 == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_1_tdata_T_58 = 8'h2 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_1_tdata_T_60 = _in_data_1_tdata_T_58 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_61 = _in_data_1_tdata_T_54 ? in_m_axis_tdata[479:448] : _in_data_1_tdata_T_60; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_62 = _in_data_1_tdata_T_50 ? in_m_axis_tdata[447:416] : _in_data_1_tdata_T_61; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_63 = _in_data_1_tdata_T_46 ? in_m_axis_tdata[415:384] : _in_data_1_tdata_T_62; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_64 = _in_data_1_tdata_T_42 ? in_m_axis_tdata[383:352] : _in_data_1_tdata_T_63; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_65 = _in_data_1_tdata_T_38 ? in_m_axis_tdata[351:320] : _in_data_1_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_66 = _in_data_1_tdata_T_34 ? in_m_axis_tdata[319:288] : _in_data_1_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_67 = _in_data_1_tdata_T_30 ? in_m_axis_tdata[287:256] : _in_data_1_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_68 = _in_data_1_tdata_T_26 ? in_m_axis_tdata[255:224] : _in_data_1_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_69 = _in_data_1_tdata_T_22 ? in_m_axis_tdata[223:192] : _in_data_1_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_70 = _in_data_1_tdata_T_18 ? in_m_axis_tdata[191:160] : _in_data_1_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_71 = _in_data_1_tdata_T_14 ? in_m_axis_tdata[159:128] : _in_data_1_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_72 = _in_data_1_tdata_T_10 ? in_m_axis_tdata[127:96] : _in_data_1_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _in_data_1_tdata_T_73 = _in_data_1_tdata_T_6 ? in_m_axis_tdata[95:64] : _in_data_1_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] in_data_1_tdata = _in_data_1_tdata_T_2 ? in_m_axis_tdata[63:32] : _in_data_1_tdata_T_73; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_61 = _in_data_1_tdata_T_54 ? in_m_axis_tkeep[14] : _in_data_1_tdata_T_58 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_62 = _in_data_1_tdata_T_50 ? in_m_axis_tkeep[13] : _in_data_1_tkeep_T_61; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_63 = _in_data_1_tdata_T_46 ? in_m_axis_tkeep[12] : _in_data_1_tkeep_T_62; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_64 = _in_data_1_tdata_T_42 ? in_m_axis_tkeep[11] : _in_data_1_tkeep_T_63; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_65 = _in_data_1_tdata_T_38 ? in_m_axis_tkeep[10] : _in_data_1_tkeep_T_64; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_66 = _in_data_1_tdata_T_34 ? in_m_axis_tkeep[9] : _in_data_1_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_67 = _in_data_1_tdata_T_30 ? in_m_axis_tkeep[8] : _in_data_1_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_68 = _in_data_1_tdata_T_26 ? in_m_axis_tkeep[7] : _in_data_1_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_69 = _in_data_1_tdata_T_22 ? in_m_axis_tkeep[6] : _in_data_1_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_70 = _in_data_1_tdata_T_18 ? in_m_axis_tkeep[5] : _in_data_1_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_71 = _in_data_1_tdata_T_14 ? in_m_axis_tkeep[4] : _in_data_1_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_72 = _in_data_1_tdata_T_10 ? in_m_axis_tkeep[3] : _in_data_1_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _in_data_1_tkeep_T_73 = _in_data_1_tdata_T_6 ? in_m_axis_tkeep[2] : _in_data_1_tkeep_T_72; // @[Mux.scala 98:16]
  wire  in_data_1_tkeep = _in_data_1_tdata_T_2 ? in_m_axis_tkeep[1] : _in_data_1_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _in_data_2_tdata_T_2 = 8'h3 == in_count_2; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_6 = 8'h3 == in_count_3; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_10 = 8'h3 == in_count_4; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_14 = 8'h3 == in_count_5; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_18 = 8'h3 == in_count_6; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_22 = 8'h3 == in_count_7; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_26 = 8'h3 == in_count_8; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_30 = 8'h3 == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_34 = 8'h3 == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_38 = 8'h3 == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_42 = 8'h3 == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_46 = 8'h3 == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_50 = 8'h3 == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_2_tdata_T_54 = 8'h3 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_2_tdata_T_56 = _in_data_2_tdata_T_54 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_57 = _in_data_2_tdata_T_50 ? in_m_axis_tdata[479:448] : _in_data_2_tdata_T_56; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_58 = _in_data_2_tdata_T_46 ? in_m_axis_tdata[447:416] : _in_data_2_tdata_T_57; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_59 = _in_data_2_tdata_T_42 ? in_m_axis_tdata[415:384] : _in_data_2_tdata_T_58; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_60 = _in_data_2_tdata_T_38 ? in_m_axis_tdata[383:352] : _in_data_2_tdata_T_59; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_61 = _in_data_2_tdata_T_34 ? in_m_axis_tdata[351:320] : _in_data_2_tdata_T_60; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_62 = _in_data_2_tdata_T_30 ? in_m_axis_tdata[319:288] : _in_data_2_tdata_T_61; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_63 = _in_data_2_tdata_T_26 ? in_m_axis_tdata[287:256] : _in_data_2_tdata_T_62; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_64 = _in_data_2_tdata_T_22 ? in_m_axis_tdata[255:224] : _in_data_2_tdata_T_63; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_65 = _in_data_2_tdata_T_18 ? in_m_axis_tdata[223:192] : _in_data_2_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_66 = _in_data_2_tdata_T_14 ? in_m_axis_tdata[191:160] : _in_data_2_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_67 = _in_data_2_tdata_T_10 ? in_m_axis_tdata[159:128] : _in_data_2_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _in_data_2_tdata_T_68 = _in_data_2_tdata_T_6 ? in_m_axis_tdata[127:96] : _in_data_2_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] in_data_2_tdata = _in_data_2_tdata_T_2 ? in_m_axis_tdata[95:64] : _in_data_2_tdata_T_68; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_57 = _in_data_2_tdata_T_50 ? in_m_axis_tkeep[14] : _in_data_2_tdata_T_54 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_58 = _in_data_2_tdata_T_46 ? in_m_axis_tkeep[13] : _in_data_2_tkeep_T_57; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_59 = _in_data_2_tdata_T_42 ? in_m_axis_tkeep[12] : _in_data_2_tkeep_T_58; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_60 = _in_data_2_tdata_T_38 ? in_m_axis_tkeep[11] : _in_data_2_tkeep_T_59; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_61 = _in_data_2_tdata_T_34 ? in_m_axis_tkeep[10] : _in_data_2_tkeep_T_60; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_62 = _in_data_2_tdata_T_30 ? in_m_axis_tkeep[9] : _in_data_2_tkeep_T_61; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_63 = _in_data_2_tdata_T_26 ? in_m_axis_tkeep[8] : _in_data_2_tkeep_T_62; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_64 = _in_data_2_tdata_T_22 ? in_m_axis_tkeep[7] : _in_data_2_tkeep_T_63; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_65 = _in_data_2_tdata_T_18 ? in_m_axis_tkeep[6] : _in_data_2_tkeep_T_64; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_66 = _in_data_2_tdata_T_14 ? in_m_axis_tkeep[5] : _in_data_2_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_67 = _in_data_2_tdata_T_10 ? in_m_axis_tkeep[4] : _in_data_2_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _in_data_2_tkeep_T_68 = _in_data_2_tdata_T_6 ? in_m_axis_tkeep[3] : _in_data_2_tkeep_T_67; // @[Mux.scala 98:16]
  wire  in_data_2_tkeep = _in_data_2_tdata_T_2 ? in_m_axis_tkeep[2] : _in_data_2_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _in_data_3_tdata_T_2 = 8'h4 == in_count_3; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_6 = 8'h4 == in_count_4; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_10 = 8'h4 == in_count_5; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_14 = 8'h4 == in_count_6; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_18 = 8'h4 == in_count_7; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_22 = 8'h4 == in_count_8; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_26 = 8'h4 == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_30 = 8'h4 == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_34 = 8'h4 == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_38 = 8'h4 == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_42 = 8'h4 == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_46 = 8'h4 == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_3_tdata_T_50 = 8'h4 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_3_tdata_T_52 = _in_data_3_tdata_T_50 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_53 = _in_data_3_tdata_T_46 ? in_m_axis_tdata[479:448] : _in_data_3_tdata_T_52; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_54 = _in_data_3_tdata_T_42 ? in_m_axis_tdata[447:416] : _in_data_3_tdata_T_53; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_55 = _in_data_3_tdata_T_38 ? in_m_axis_tdata[415:384] : _in_data_3_tdata_T_54; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_56 = _in_data_3_tdata_T_34 ? in_m_axis_tdata[383:352] : _in_data_3_tdata_T_55; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_57 = _in_data_3_tdata_T_30 ? in_m_axis_tdata[351:320] : _in_data_3_tdata_T_56; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_58 = _in_data_3_tdata_T_26 ? in_m_axis_tdata[319:288] : _in_data_3_tdata_T_57; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_59 = _in_data_3_tdata_T_22 ? in_m_axis_tdata[287:256] : _in_data_3_tdata_T_58; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_60 = _in_data_3_tdata_T_18 ? in_m_axis_tdata[255:224] : _in_data_3_tdata_T_59; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_61 = _in_data_3_tdata_T_14 ? in_m_axis_tdata[223:192] : _in_data_3_tdata_T_60; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_62 = _in_data_3_tdata_T_10 ? in_m_axis_tdata[191:160] : _in_data_3_tdata_T_61; // @[Mux.scala 98:16]
  wire [31:0] _in_data_3_tdata_T_63 = _in_data_3_tdata_T_6 ? in_m_axis_tdata[159:128] : _in_data_3_tdata_T_62; // @[Mux.scala 98:16]
  wire [31:0] in_data_3_tdata = _in_data_3_tdata_T_2 ? in_m_axis_tdata[127:96] : _in_data_3_tdata_T_63; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_53 = _in_data_3_tdata_T_46 ? in_m_axis_tkeep[14] : _in_data_3_tdata_T_50 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_54 = _in_data_3_tdata_T_42 ? in_m_axis_tkeep[13] : _in_data_3_tkeep_T_53; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_55 = _in_data_3_tdata_T_38 ? in_m_axis_tkeep[12] : _in_data_3_tkeep_T_54; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_56 = _in_data_3_tdata_T_34 ? in_m_axis_tkeep[11] : _in_data_3_tkeep_T_55; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_57 = _in_data_3_tdata_T_30 ? in_m_axis_tkeep[10] : _in_data_3_tkeep_T_56; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_58 = _in_data_3_tdata_T_26 ? in_m_axis_tkeep[9] : _in_data_3_tkeep_T_57; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_59 = _in_data_3_tdata_T_22 ? in_m_axis_tkeep[8] : _in_data_3_tkeep_T_58; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_60 = _in_data_3_tdata_T_18 ? in_m_axis_tkeep[7] : _in_data_3_tkeep_T_59; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_61 = _in_data_3_tdata_T_14 ? in_m_axis_tkeep[6] : _in_data_3_tkeep_T_60; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_62 = _in_data_3_tdata_T_10 ? in_m_axis_tkeep[5] : _in_data_3_tkeep_T_61; // @[Mux.scala 98:16]
  wire  _in_data_3_tkeep_T_63 = _in_data_3_tdata_T_6 ? in_m_axis_tkeep[4] : _in_data_3_tkeep_T_62; // @[Mux.scala 98:16]
  wire  in_data_3_tkeep = _in_data_3_tdata_T_2 ? in_m_axis_tkeep[3] : _in_data_3_tkeep_T_63; // @[Mux.scala 98:16]
  wire  _in_data_4_tdata_T_2 = 8'h5 == in_count_4; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_6 = 8'h5 == in_count_5; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_10 = 8'h5 == in_count_6; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_14 = 8'h5 == in_count_7; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_18 = 8'h5 == in_count_8; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_22 = 8'h5 == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_26 = 8'h5 == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_30 = 8'h5 == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_34 = 8'h5 == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_38 = 8'h5 == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_42 = 8'h5 == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_4_tdata_T_46 = 8'h5 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_4_tdata_T_48 = _in_data_4_tdata_T_46 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_49 = _in_data_4_tdata_T_42 ? in_m_axis_tdata[479:448] : _in_data_4_tdata_T_48; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_50 = _in_data_4_tdata_T_38 ? in_m_axis_tdata[447:416] : _in_data_4_tdata_T_49; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_51 = _in_data_4_tdata_T_34 ? in_m_axis_tdata[415:384] : _in_data_4_tdata_T_50; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_52 = _in_data_4_tdata_T_30 ? in_m_axis_tdata[383:352] : _in_data_4_tdata_T_51; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_53 = _in_data_4_tdata_T_26 ? in_m_axis_tdata[351:320] : _in_data_4_tdata_T_52; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_54 = _in_data_4_tdata_T_22 ? in_m_axis_tdata[319:288] : _in_data_4_tdata_T_53; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_55 = _in_data_4_tdata_T_18 ? in_m_axis_tdata[287:256] : _in_data_4_tdata_T_54; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_56 = _in_data_4_tdata_T_14 ? in_m_axis_tdata[255:224] : _in_data_4_tdata_T_55; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_57 = _in_data_4_tdata_T_10 ? in_m_axis_tdata[223:192] : _in_data_4_tdata_T_56; // @[Mux.scala 98:16]
  wire [31:0] _in_data_4_tdata_T_58 = _in_data_4_tdata_T_6 ? in_m_axis_tdata[191:160] : _in_data_4_tdata_T_57; // @[Mux.scala 98:16]
  wire [31:0] in_data_4_tdata = _in_data_4_tdata_T_2 ? in_m_axis_tdata[159:128] : _in_data_4_tdata_T_58; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_49 = _in_data_4_tdata_T_42 ? in_m_axis_tkeep[14] : _in_data_4_tdata_T_46 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_50 = _in_data_4_tdata_T_38 ? in_m_axis_tkeep[13] : _in_data_4_tkeep_T_49; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_51 = _in_data_4_tdata_T_34 ? in_m_axis_tkeep[12] : _in_data_4_tkeep_T_50; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_52 = _in_data_4_tdata_T_30 ? in_m_axis_tkeep[11] : _in_data_4_tkeep_T_51; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_53 = _in_data_4_tdata_T_26 ? in_m_axis_tkeep[10] : _in_data_4_tkeep_T_52; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_54 = _in_data_4_tdata_T_22 ? in_m_axis_tkeep[9] : _in_data_4_tkeep_T_53; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_55 = _in_data_4_tdata_T_18 ? in_m_axis_tkeep[8] : _in_data_4_tkeep_T_54; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_56 = _in_data_4_tdata_T_14 ? in_m_axis_tkeep[7] : _in_data_4_tkeep_T_55; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_57 = _in_data_4_tdata_T_10 ? in_m_axis_tkeep[6] : _in_data_4_tkeep_T_56; // @[Mux.scala 98:16]
  wire  _in_data_4_tkeep_T_58 = _in_data_4_tdata_T_6 ? in_m_axis_tkeep[5] : _in_data_4_tkeep_T_57; // @[Mux.scala 98:16]
  wire  in_data_4_tkeep = _in_data_4_tdata_T_2 ? in_m_axis_tkeep[4] : _in_data_4_tkeep_T_58; // @[Mux.scala 98:16]
  wire  _in_data_5_tdata_T_2 = 8'h6 == in_count_5; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_6 = 8'h6 == in_count_6; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_10 = 8'h6 == in_count_7; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_14 = 8'h6 == in_count_8; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_18 = 8'h6 == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_22 = 8'h6 == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_26 = 8'h6 == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_30 = 8'h6 == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_34 = 8'h6 == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_38 = 8'h6 == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_5_tdata_T_42 = 8'h6 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_5_tdata_T_44 = _in_data_5_tdata_T_42 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_5_tdata_T_45 = _in_data_5_tdata_T_38 ? in_m_axis_tdata[479:448] : _in_data_5_tdata_T_44; // @[Mux.scala 98:16]
  wire [31:0] _in_data_5_tdata_T_46 = _in_data_5_tdata_T_34 ? in_m_axis_tdata[447:416] : _in_data_5_tdata_T_45; // @[Mux.scala 98:16]
  wire [31:0] _in_data_5_tdata_T_47 = _in_data_5_tdata_T_30 ? in_m_axis_tdata[415:384] : _in_data_5_tdata_T_46; // @[Mux.scala 98:16]
  wire [31:0] _in_data_5_tdata_T_48 = _in_data_5_tdata_T_26 ? in_m_axis_tdata[383:352] : _in_data_5_tdata_T_47; // @[Mux.scala 98:16]
  wire [31:0] _in_data_5_tdata_T_49 = _in_data_5_tdata_T_22 ? in_m_axis_tdata[351:320] : _in_data_5_tdata_T_48; // @[Mux.scala 98:16]
  wire [31:0] _in_data_5_tdata_T_50 = _in_data_5_tdata_T_18 ? in_m_axis_tdata[319:288] : _in_data_5_tdata_T_49; // @[Mux.scala 98:16]
  wire [31:0] _in_data_5_tdata_T_51 = _in_data_5_tdata_T_14 ? in_m_axis_tdata[287:256] : _in_data_5_tdata_T_50; // @[Mux.scala 98:16]
  wire [31:0] _in_data_5_tdata_T_52 = _in_data_5_tdata_T_10 ? in_m_axis_tdata[255:224] : _in_data_5_tdata_T_51; // @[Mux.scala 98:16]
  wire [31:0] _in_data_5_tdata_T_53 = _in_data_5_tdata_T_6 ? in_m_axis_tdata[223:192] : _in_data_5_tdata_T_52; // @[Mux.scala 98:16]
  wire [31:0] in_data_5_tdata = _in_data_5_tdata_T_2 ? in_m_axis_tdata[191:160] : _in_data_5_tdata_T_53; // @[Mux.scala 98:16]
  wire  _in_data_5_tkeep_T_45 = _in_data_5_tdata_T_38 ? in_m_axis_tkeep[14] : _in_data_5_tdata_T_42 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_5_tkeep_T_46 = _in_data_5_tdata_T_34 ? in_m_axis_tkeep[13] : _in_data_5_tkeep_T_45; // @[Mux.scala 98:16]
  wire  _in_data_5_tkeep_T_47 = _in_data_5_tdata_T_30 ? in_m_axis_tkeep[12] : _in_data_5_tkeep_T_46; // @[Mux.scala 98:16]
  wire  _in_data_5_tkeep_T_48 = _in_data_5_tdata_T_26 ? in_m_axis_tkeep[11] : _in_data_5_tkeep_T_47; // @[Mux.scala 98:16]
  wire  _in_data_5_tkeep_T_49 = _in_data_5_tdata_T_22 ? in_m_axis_tkeep[10] : _in_data_5_tkeep_T_48; // @[Mux.scala 98:16]
  wire  _in_data_5_tkeep_T_50 = _in_data_5_tdata_T_18 ? in_m_axis_tkeep[9] : _in_data_5_tkeep_T_49; // @[Mux.scala 98:16]
  wire  _in_data_5_tkeep_T_51 = _in_data_5_tdata_T_14 ? in_m_axis_tkeep[8] : _in_data_5_tkeep_T_50; // @[Mux.scala 98:16]
  wire  _in_data_5_tkeep_T_52 = _in_data_5_tdata_T_10 ? in_m_axis_tkeep[7] : _in_data_5_tkeep_T_51; // @[Mux.scala 98:16]
  wire  _in_data_5_tkeep_T_53 = _in_data_5_tdata_T_6 ? in_m_axis_tkeep[6] : _in_data_5_tkeep_T_52; // @[Mux.scala 98:16]
  wire  in_data_5_tkeep = _in_data_5_tdata_T_2 ? in_m_axis_tkeep[5] : _in_data_5_tkeep_T_53; // @[Mux.scala 98:16]
  wire  _in_data_6_tdata_T_2 = 8'h7 == in_count_6; // @[bfs_remote.scala 35:37]
  wire  _in_data_6_tdata_T_6 = 8'h7 == in_count_7; // @[bfs_remote.scala 35:37]
  wire  _in_data_6_tdata_T_10 = 8'h7 == in_count_8; // @[bfs_remote.scala 35:37]
  wire  _in_data_6_tdata_T_14 = 8'h7 == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_6_tdata_T_18 = 8'h7 == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_6_tdata_T_22 = 8'h7 == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_6_tdata_T_26 = 8'h7 == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_6_tdata_T_30 = 8'h7 == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_6_tdata_T_34 = 8'h7 == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_6_tdata_T_38 = 8'h7 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_6_tdata_T_40 = _in_data_6_tdata_T_38 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_6_tdata_T_41 = _in_data_6_tdata_T_34 ? in_m_axis_tdata[479:448] : _in_data_6_tdata_T_40; // @[Mux.scala 98:16]
  wire [31:0] _in_data_6_tdata_T_42 = _in_data_6_tdata_T_30 ? in_m_axis_tdata[447:416] : _in_data_6_tdata_T_41; // @[Mux.scala 98:16]
  wire [31:0] _in_data_6_tdata_T_43 = _in_data_6_tdata_T_26 ? in_m_axis_tdata[415:384] : _in_data_6_tdata_T_42; // @[Mux.scala 98:16]
  wire [31:0] _in_data_6_tdata_T_44 = _in_data_6_tdata_T_22 ? in_m_axis_tdata[383:352] : _in_data_6_tdata_T_43; // @[Mux.scala 98:16]
  wire [31:0] _in_data_6_tdata_T_45 = _in_data_6_tdata_T_18 ? in_m_axis_tdata[351:320] : _in_data_6_tdata_T_44; // @[Mux.scala 98:16]
  wire [31:0] _in_data_6_tdata_T_46 = _in_data_6_tdata_T_14 ? in_m_axis_tdata[319:288] : _in_data_6_tdata_T_45; // @[Mux.scala 98:16]
  wire [31:0] _in_data_6_tdata_T_47 = _in_data_6_tdata_T_10 ? in_m_axis_tdata[287:256] : _in_data_6_tdata_T_46; // @[Mux.scala 98:16]
  wire [31:0] _in_data_6_tdata_T_48 = _in_data_6_tdata_T_6 ? in_m_axis_tdata[255:224] : _in_data_6_tdata_T_47; // @[Mux.scala 98:16]
  wire [31:0] in_data_6_tdata = _in_data_6_tdata_T_2 ? in_m_axis_tdata[223:192] : _in_data_6_tdata_T_48; // @[Mux.scala 98:16]
  wire  _in_data_6_tkeep_T_41 = _in_data_6_tdata_T_34 ? in_m_axis_tkeep[14] : _in_data_6_tdata_T_38 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_6_tkeep_T_42 = _in_data_6_tdata_T_30 ? in_m_axis_tkeep[13] : _in_data_6_tkeep_T_41; // @[Mux.scala 98:16]
  wire  _in_data_6_tkeep_T_43 = _in_data_6_tdata_T_26 ? in_m_axis_tkeep[12] : _in_data_6_tkeep_T_42; // @[Mux.scala 98:16]
  wire  _in_data_6_tkeep_T_44 = _in_data_6_tdata_T_22 ? in_m_axis_tkeep[11] : _in_data_6_tkeep_T_43; // @[Mux.scala 98:16]
  wire  _in_data_6_tkeep_T_45 = _in_data_6_tdata_T_18 ? in_m_axis_tkeep[10] : _in_data_6_tkeep_T_44; // @[Mux.scala 98:16]
  wire  _in_data_6_tkeep_T_46 = _in_data_6_tdata_T_14 ? in_m_axis_tkeep[9] : _in_data_6_tkeep_T_45; // @[Mux.scala 98:16]
  wire  _in_data_6_tkeep_T_47 = _in_data_6_tdata_T_10 ? in_m_axis_tkeep[8] : _in_data_6_tkeep_T_46; // @[Mux.scala 98:16]
  wire  _in_data_6_tkeep_T_48 = _in_data_6_tdata_T_6 ? in_m_axis_tkeep[7] : _in_data_6_tkeep_T_47; // @[Mux.scala 98:16]
  wire  in_data_6_tkeep = _in_data_6_tdata_T_2 ? in_m_axis_tkeep[6] : _in_data_6_tkeep_T_48; // @[Mux.scala 98:16]
  wire  _in_data_7_tdata_T_2 = 8'h8 == in_count_7; // @[bfs_remote.scala 35:37]
  wire  _in_data_7_tdata_T_6 = 8'h8 == in_count_8; // @[bfs_remote.scala 35:37]
  wire  _in_data_7_tdata_T_10 = 8'h8 == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_7_tdata_T_14 = 8'h8 == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_7_tdata_T_18 = 8'h8 == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_7_tdata_T_22 = 8'h8 == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_7_tdata_T_26 = 8'h8 == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_7_tdata_T_30 = 8'h8 == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_7_tdata_T_34 = 8'h8 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_7_tdata_T_36 = _in_data_7_tdata_T_34 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_7_tdata_T_37 = _in_data_7_tdata_T_30 ? in_m_axis_tdata[479:448] : _in_data_7_tdata_T_36; // @[Mux.scala 98:16]
  wire [31:0] _in_data_7_tdata_T_38 = _in_data_7_tdata_T_26 ? in_m_axis_tdata[447:416] : _in_data_7_tdata_T_37; // @[Mux.scala 98:16]
  wire [31:0] _in_data_7_tdata_T_39 = _in_data_7_tdata_T_22 ? in_m_axis_tdata[415:384] : _in_data_7_tdata_T_38; // @[Mux.scala 98:16]
  wire [31:0] _in_data_7_tdata_T_40 = _in_data_7_tdata_T_18 ? in_m_axis_tdata[383:352] : _in_data_7_tdata_T_39; // @[Mux.scala 98:16]
  wire [31:0] _in_data_7_tdata_T_41 = _in_data_7_tdata_T_14 ? in_m_axis_tdata[351:320] : _in_data_7_tdata_T_40; // @[Mux.scala 98:16]
  wire [31:0] _in_data_7_tdata_T_42 = _in_data_7_tdata_T_10 ? in_m_axis_tdata[319:288] : _in_data_7_tdata_T_41; // @[Mux.scala 98:16]
  wire [31:0] _in_data_7_tdata_T_43 = _in_data_7_tdata_T_6 ? in_m_axis_tdata[287:256] : _in_data_7_tdata_T_42; // @[Mux.scala 98:16]
  wire [31:0] in_data_7_tdata = _in_data_7_tdata_T_2 ? in_m_axis_tdata[255:224] : _in_data_7_tdata_T_43; // @[Mux.scala 98:16]
  wire  _in_data_7_tkeep_T_37 = _in_data_7_tdata_T_30 ? in_m_axis_tkeep[14] : _in_data_7_tdata_T_34 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_7_tkeep_T_38 = _in_data_7_tdata_T_26 ? in_m_axis_tkeep[13] : _in_data_7_tkeep_T_37; // @[Mux.scala 98:16]
  wire  _in_data_7_tkeep_T_39 = _in_data_7_tdata_T_22 ? in_m_axis_tkeep[12] : _in_data_7_tkeep_T_38; // @[Mux.scala 98:16]
  wire  _in_data_7_tkeep_T_40 = _in_data_7_tdata_T_18 ? in_m_axis_tkeep[11] : _in_data_7_tkeep_T_39; // @[Mux.scala 98:16]
  wire  _in_data_7_tkeep_T_41 = _in_data_7_tdata_T_14 ? in_m_axis_tkeep[10] : _in_data_7_tkeep_T_40; // @[Mux.scala 98:16]
  wire  _in_data_7_tkeep_T_42 = _in_data_7_tdata_T_10 ? in_m_axis_tkeep[9] : _in_data_7_tkeep_T_41; // @[Mux.scala 98:16]
  wire  _in_data_7_tkeep_T_43 = _in_data_7_tdata_T_6 ? in_m_axis_tkeep[8] : _in_data_7_tkeep_T_42; // @[Mux.scala 98:16]
  wire  in_data_7_tkeep = _in_data_7_tdata_T_2 ? in_m_axis_tkeep[7] : _in_data_7_tkeep_T_43; // @[Mux.scala 98:16]
  wire  _in_data_8_tdata_T_2 = 8'h9 == in_count_8; // @[bfs_remote.scala 35:37]
  wire  _in_data_8_tdata_T_6 = 8'h9 == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_8_tdata_T_10 = 8'h9 == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_8_tdata_T_14 = 8'h9 == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_8_tdata_T_18 = 8'h9 == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_8_tdata_T_22 = 8'h9 == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_8_tdata_T_26 = 8'h9 == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_8_tdata_T_30 = 8'h9 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_8_tdata_T_32 = _in_data_8_tdata_T_30 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_8_tdata_T_33 = _in_data_8_tdata_T_26 ? in_m_axis_tdata[479:448] : _in_data_8_tdata_T_32; // @[Mux.scala 98:16]
  wire [31:0] _in_data_8_tdata_T_34 = _in_data_8_tdata_T_22 ? in_m_axis_tdata[447:416] : _in_data_8_tdata_T_33; // @[Mux.scala 98:16]
  wire [31:0] _in_data_8_tdata_T_35 = _in_data_8_tdata_T_18 ? in_m_axis_tdata[415:384] : _in_data_8_tdata_T_34; // @[Mux.scala 98:16]
  wire [31:0] _in_data_8_tdata_T_36 = _in_data_8_tdata_T_14 ? in_m_axis_tdata[383:352] : _in_data_8_tdata_T_35; // @[Mux.scala 98:16]
  wire [31:0] _in_data_8_tdata_T_37 = _in_data_8_tdata_T_10 ? in_m_axis_tdata[351:320] : _in_data_8_tdata_T_36; // @[Mux.scala 98:16]
  wire [31:0] _in_data_8_tdata_T_38 = _in_data_8_tdata_T_6 ? in_m_axis_tdata[319:288] : _in_data_8_tdata_T_37; // @[Mux.scala 98:16]
  wire [31:0] in_data_8_tdata = _in_data_8_tdata_T_2 ? in_m_axis_tdata[287:256] : _in_data_8_tdata_T_38; // @[Mux.scala 98:16]
  wire  _in_data_8_tkeep_T_33 = _in_data_8_tdata_T_26 ? in_m_axis_tkeep[14] : _in_data_8_tdata_T_30 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_8_tkeep_T_34 = _in_data_8_tdata_T_22 ? in_m_axis_tkeep[13] : _in_data_8_tkeep_T_33; // @[Mux.scala 98:16]
  wire  _in_data_8_tkeep_T_35 = _in_data_8_tdata_T_18 ? in_m_axis_tkeep[12] : _in_data_8_tkeep_T_34; // @[Mux.scala 98:16]
  wire  _in_data_8_tkeep_T_36 = _in_data_8_tdata_T_14 ? in_m_axis_tkeep[11] : _in_data_8_tkeep_T_35; // @[Mux.scala 98:16]
  wire  _in_data_8_tkeep_T_37 = _in_data_8_tdata_T_10 ? in_m_axis_tkeep[10] : _in_data_8_tkeep_T_36; // @[Mux.scala 98:16]
  wire  _in_data_8_tkeep_T_38 = _in_data_8_tdata_T_6 ? in_m_axis_tkeep[9] : _in_data_8_tkeep_T_37; // @[Mux.scala 98:16]
  wire  in_data_8_tkeep = _in_data_8_tdata_T_2 ? in_m_axis_tkeep[8] : _in_data_8_tkeep_T_38; // @[Mux.scala 98:16]
  wire  _in_data_9_tdata_T_2 = 8'ha == in_count_9; // @[bfs_remote.scala 35:37]
  wire  _in_data_9_tdata_T_6 = 8'ha == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_9_tdata_T_10 = 8'ha == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_9_tdata_T_14 = 8'ha == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_9_tdata_T_18 = 8'ha == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_9_tdata_T_22 = 8'ha == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_9_tdata_T_26 = 8'ha == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_9_tdata_T_28 = _in_data_9_tdata_T_26 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_9_tdata_T_29 = _in_data_9_tdata_T_22 ? in_m_axis_tdata[479:448] : _in_data_9_tdata_T_28; // @[Mux.scala 98:16]
  wire [31:0] _in_data_9_tdata_T_30 = _in_data_9_tdata_T_18 ? in_m_axis_tdata[447:416] : _in_data_9_tdata_T_29; // @[Mux.scala 98:16]
  wire [31:0] _in_data_9_tdata_T_31 = _in_data_9_tdata_T_14 ? in_m_axis_tdata[415:384] : _in_data_9_tdata_T_30; // @[Mux.scala 98:16]
  wire [31:0] _in_data_9_tdata_T_32 = _in_data_9_tdata_T_10 ? in_m_axis_tdata[383:352] : _in_data_9_tdata_T_31; // @[Mux.scala 98:16]
  wire [31:0] _in_data_9_tdata_T_33 = _in_data_9_tdata_T_6 ? in_m_axis_tdata[351:320] : _in_data_9_tdata_T_32; // @[Mux.scala 98:16]
  wire [31:0] in_data_9_tdata = _in_data_9_tdata_T_2 ? in_m_axis_tdata[319:288] : _in_data_9_tdata_T_33; // @[Mux.scala 98:16]
  wire  _in_data_9_tkeep_T_29 = _in_data_9_tdata_T_22 ? in_m_axis_tkeep[14] : _in_data_9_tdata_T_26 & in_m_axis_tkeep[15
    ]; // @[Mux.scala 98:16]
  wire  _in_data_9_tkeep_T_30 = _in_data_9_tdata_T_18 ? in_m_axis_tkeep[13] : _in_data_9_tkeep_T_29; // @[Mux.scala 98:16]
  wire  _in_data_9_tkeep_T_31 = _in_data_9_tdata_T_14 ? in_m_axis_tkeep[12] : _in_data_9_tkeep_T_30; // @[Mux.scala 98:16]
  wire  _in_data_9_tkeep_T_32 = _in_data_9_tdata_T_10 ? in_m_axis_tkeep[11] : _in_data_9_tkeep_T_31; // @[Mux.scala 98:16]
  wire  _in_data_9_tkeep_T_33 = _in_data_9_tdata_T_6 ? in_m_axis_tkeep[10] : _in_data_9_tkeep_T_32; // @[Mux.scala 98:16]
  wire  in_data_9_tkeep = _in_data_9_tdata_T_2 ? in_m_axis_tkeep[9] : _in_data_9_tkeep_T_33; // @[Mux.scala 98:16]
  wire  _in_data_10_tdata_T_2 = 8'hb == in_count_10; // @[bfs_remote.scala 35:37]
  wire  _in_data_10_tdata_T_6 = 8'hb == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_10_tdata_T_10 = 8'hb == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_10_tdata_T_14 = 8'hb == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_10_tdata_T_18 = 8'hb == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_10_tdata_T_22 = 8'hb == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_10_tdata_T_24 = _in_data_10_tdata_T_22 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_10_tdata_T_25 = _in_data_10_tdata_T_18 ? in_m_axis_tdata[479:448] : _in_data_10_tdata_T_24; // @[Mux.scala 98:16]
  wire [31:0] _in_data_10_tdata_T_26 = _in_data_10_tdata_T_14 ? in_m_axis_tdata[447:416] : _in_data_10_tdata_T_25; // @[Mux.scala 98:16]
  wire [31:0] _in_data_10_tdata_T_27 = _in_data_10_tdata_T_10 ? in_m_axis_tdata[415:384] : _in_data_10_tdata_T_26; // @[Mux.scala 98:16]
  wire [31:0] _in_data_10_tdata_T_28 = _in_data_10_tdata_T_6 ? in_m_axis_tdata[383:352] : _in_data_10_tdata_T_27; // @[Mux.scala 98:16]
  wire [31:0] in_data_10_tdata = _in_data_10_tdata_T_2 ? in_m_axis_tdata[351:320] : _in_data_10_tdata_T_28; // @[Mux.scala 98:16]
  wire  _in_data_10_tkeep_T_25 = _in_data_10_tdata_T_18 ? in_m_axis_tkeep[14] : _in_data_10_tdata_T_22 & in_m_axis_tkeep
    [15]; // @[Mux.scala 98:16]
  wire  _in_data_10_tkeep_T_26 = _in_data_10_tdata_T_14 ? in_m_axis_tkeep[13] : _in_data_10_tkeep_T_25; // @[Mux.scala 98:16]
  wire  _in_data_10_tkeep_T_27 = _in_data_10_tdata_T_10 ? in_m_axis_tkeep[12] : _in_data_10_tkeep_T_26; // @[Mux.scala 98:16]
  wire  _in_data_10_tkeep_T_28 = _in_data_10_tdata_T_6 ? in_m_axis_tkeep[11] : _in_data_10_tkeep_T_27; // @[Mux.scala 98:16]
  wire  in_data_10_tkeep = _in_data_10_tdata_T_2 ? in_m_axis_tkeep[10] : _in_data_10_tkeep_T_28; // @[Mux.scala 98:16]
  wire  _in_data_11_tdata_T_2 = 8'hc == in_count_11; // @[bfs_remote.scala 35:37]
  wire  _in_data_11_tdata_T_6 = 8'hc == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_11_tdata_T_10 = 8'hc == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_11_tdata_T_14 = 8'hc == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_11_tdata_T_18 = 8'hc == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_11_tdata_T_20 = _in_data_11_tdata_T_18 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_11_tdata_T_21 = _in_data_11_tdata_T_14 ? in_m_axis_tdata[479:448] : _in_data_11_tdata_T_20; // @[Mux.scala 98:16]
  wire [31:0] _in_data_11_tdata_T_22 = _in_data_11_tdata_T_10 ? in_m_axis_tdata[447:416] : _in_data_11_tdata_T_21; // @[Mux.scala 98:16]
  wire [31:0] _in_data_11_tdata_T_23 = _in_data_11_tdata_T_6 ? in_m_axis_tdata[415:384] : _in_data_11_tdata_T_22; // @[Mux.scala 98:16]
  wire [31:0] in_data_11_tdata = _in_data_11_tdata_T_2 ? in_m_axis_tdata[383:352] : _in_data_11_tdata_T_23; // @[Mux.scala 98:16]
  wire  _in_data_11_tkeep_T_21 = _in_data_11_tdata_T_14 ? in_m_axis_tkeep[14] : _in_data_11_tdata_T_18 & in_m_axis_tkeep
    [15]; // @[Mux.scala 98:16]
  wire  _in_data_11_tkeep_T_22 = _in_data_11_tdata_T_10 ? in_m_axis_tkeep[13] : _in_data_11_tkeep_T_21; // @[Mux.scala 98:16]
  wire  _in_data_11_tkeep_T_23 = _in_data_11_tdata_T_6 ? in_m_axis_tkeep[12] : _in_data_11_tkeep_T_22; // @[Mux.scala 98:16]
  wire  in_data_11_tkeep = _in_data_11_tdata_T_2 ? in_m_axis_tkeep[11] : _in_data_11_tkeep_T_23; // @[Mux.scala 98:16]
  wire  _in_data_12_tdata_T_2 = 8'hd == in_count_12; // @[bfs_remote.scala 35:37]
  wire  _in_data_12_tdata_T_6 = 8'hd == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_12_tdata_T_10 = 8'hd == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_12_tdata_T_14 = 8'hd == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_12_tdata_T_16 = _in_data_12_tdata_T_14 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_12_tdata_T_17 = _in_data_12_tdata_T_10 ? in_m_axis_tdata[479:448] : _in_data_12_tdata_T_16; // @[Mux.scala 98:16]
  wire [31:0] _in_data_12_tdata_T_18 = _in_data_12_tdata_T_6 ? in_m_axis_tdata[447:416] : _in_data_12_tdata_T_17; // @[Mux.scala 98:16]
  wire [31:0] in_data_12_tdata = _in_data_12_tdata_T_2 ? in_m_axis_tdata[415:384] : _in_data_12_tdata_T_18; // @[Mux.scala 98:16]
  wire  _in_data_12_tkeep_T_17 = _in_data_12_tdata_T_10 ? in_m_axis_tkeep[14] : _in_data_12_tdata_T_14 & in_m_axis_tkeep
    [15]; // @[Mux.scala 98:16]
  wire  _in_data_12_tkeep_T_18 = _in_data_12_tdata_T_6 ? in_m_axis_tkeep[13] : _in_data_12_tkeep_T_17; // @[Mux.scala 98:16]
  wire  in_data_12_tkeep = _in_data_12_tdata_T_2 ? in_m_axis_tkeep[12] : _in_data_12_tkeep_T_18; // @[Mux.scala 98:16]
  wire  _in_data_13_tdata_T_2 = 8'he == in_count_13; // @[bfs_remote.scala 35:37]
  wire  _in_data_13_tdata_T_6 = 8'he == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_13_tdata_T_10 = 8'he == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_13_tdata_T_12 = _in_data_13_tdata_T_10 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _in_data_13_tdata_T_13 = _in_data_13_tdata_T_6 ? in_m_axis_tdata[479:448] : _in_data_13_tdata_T_12; // @[Mux.scala 98:16]
  wire [31:0] in_data_13_tdata = _in_data_13_tdata_T_2 ? in_m_axis_tdata[447:416] : _in_data_13_tdata_T_13; // @[Mux.scala 98:16]
  wire  _in_data_13_tkeep_T_13 = _in_data_13_tdata_T_6 ? in_m_axis_tkeep[14] : _in_data_13_tdata_T_10 & in_m_axis_tkeep[
    15]; // @[Mux.scala 98:16]
  wire  in_data_13_tkeep = _in_data_13_tdata_T_2 ? in_m_axis_tkeep[13] : _in_data_13_tkeep_T_13; // @[Mux.scala 98:16]
  wire  _in_data_14_tdata_T_2 = 8'hf == in_count_14; // @[bfs_remote.scala 35:37]
  wire  _in_data_14_tdata_T_6 = 8'hf == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] _in_data_14_tdata_T_8 = _in_data_14_tdata_T_6 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] in_data_14_tdata = _in_data_14_tdata_T_2 ? in_m_axis_tdata[479:448] : _in_data_14_tdata_T_8; // @[Mux.scala 98:16]
  wire  in_data_14_tkeep = _in_data_14_tdata_T_2 ? in_m_axis_tkeep[14] : _in_data_14_tdata_T_6 & in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _in_data_15_tdata_T_2 = 8'h10 == in_count_15; // @[bfs_remote.scala 35:37]
  wire [31:0] in_data_15_tdata = _in_data_15_tdata_T_2 ? in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire  in_data_15_tkeep = _in_data_15_tdata_T_2 & in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire [7:0] sorted_in_io_s_axis_tkeep_lo = {in_data_7_tkeep,in_data_6_tkeep,in_data_5_tkeep,in_data_4_tkeep,
    in_data_3_tkeep,in_data_2_tkeep,in_data_1_tkeep,in_data_0_tkeep}; // @[bfs_remote.scala 47:71]
  wire [15:0] _sorted_in_io_s_axis_tkeep_T = {in_data_15_tkeep,in_data_14_tkeep,in_data_13_tkeep,in_data_12_tkeep,
    in_data_11_tkeep,in_data_10_tkeep,in_data_9_tkeep,in_data_8_tkeep,sorted_in_io_s_axis_tkeep_lo}; // @[bfs_remote.scala 47:71]
  wire [255:0] sorted_in_io_s_axis_tdata_lo = {in_data_7_tdata,in_data_6_tdata,in_data_5_tdata,in_data_4_tdata,
    in_data_3_tdata,in_data_2_tdata,in_data_1_tdata,in_data_0_tdata}; // @[bfs_remote.scala 48:71]
  wire [255:0] sorted_in_io_s_axis_tdata_hi = {in_data_15_tdata,in_data_14_tdata,in_data_13_tdata,in_data_12_tdata,
    in_data_11_tdata,in_data_10_tdata,in_data_9_tdata,in_data_8_tdata}; // @[bfs_remote.scala 48:71]
  reg [31:0] in_count_reg; // @[bfs_remote.scala 50:29]
  reg [31:0] mid_count; // @[bfs_remote.scala 58:26]
  wire [31:0] _T_4 = 32'h0 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_0_tdata_T_3 = 32'h0 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_7 = 32'h1 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_11 = 32'h2 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_15 = 32'h3 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_19 = 32'h4 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_23 = 32'h5 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_27 = 32'h6 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_31 = 32'h7 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_35 = 32'h8 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_39 = 32'h9 == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_43 = 32'ha == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_47 = 32'hb == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_51 = 32'hc == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_55 = 32'hd == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_59 = 32'he == _T_4; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_0_tdata_T_63 = 32'hf == _T_4; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_0_tdata_T_65 = _mid_data_in_0_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_66 = _mid_data_in_0_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_0_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_67 = _mid_data_in_0_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_0_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_68 = _mid_data_in_0_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_0_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_69 = _mid_data_in_0_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_0_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_70 = _mid_data_in_0_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_0_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_71 = _mid_data_in_0_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_0_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_72 = _mid_data_in_0_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_0_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_73 = _mid_data_in_0_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_0_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_74 = _mid_data_in_0_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_0_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_75 = _mid_data_in_0_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_0_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_76 = _mid_data_in_0_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_0_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_77 = _mid_data_in_0_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_0_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_78 = _mid_data_in_0_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_0_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_79 = _mid_data_in_0_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_0_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_0_tdata_T_80 = _mid_data_in_0_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_0_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_66 = _mid_data_in_0_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_0_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_67 = _mid_data_in_0_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_0_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_68 = _mid_data_in_0_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_0_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_69 = _mid_data_in_0_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_0_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_70 = _mid_data_in_0_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_0_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_71 = _mid_data_in_0_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_0_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_72 = _mid_data_in_0_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_0_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_73 = _mid_data_in_0_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_0_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_74 = _mid_data_in_0_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_0_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_75 = _mid_data_in_0_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_0_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_76 = _mid_data_in_0_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_0_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_77 = _mid_data_in_0_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_0_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_78 = _mid_data_in_0_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_0_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_79 = _mid_data_in_0_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_0_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_0_tkeep_T_80 = _mid_data_in_0_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_0_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_1 = _T_4 < 32'h10 ? _mid_data_in_0_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_2 = _T_4 < 32'h10 & _mid_data_in_0_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_0_tdata = 32'h0 >= mid_count ? _GEN_1 : mid_m_axis_tdata[31:0]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_0_tkeep = 32'h0 >= mid_count ? _GEN_2 : mid_m_axis_tkeep[0]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_8 = 32'h1 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_1_tdata_T_3 = 32'h0 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_7 = 32'h1 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_11 = 32'h2 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_15 = 32'h3 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_19 = 32'h4 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_23 = 32'h5 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_27 = 32'h6 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_31 = 32'h7 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_35 = 32'h8 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_39 = 32'h9 == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_43 = 32'ha == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_47 = 32'hb == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_51 = 32'hc == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_55 = 32'hd == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_59 = 32'he == _T_8; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_1_tdata_T_63 = 32'hf == _T_8; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_1_tdata_T_65 = _mid_data_in_1_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_66 = _mid_data_in_1_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_1_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_67 = _mid_data_in_1_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_1_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_68 = _mid_data_in_1_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_1_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_69 = _mid_data_in_1_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_1_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_70 = _mid_data_in_1_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_1_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_71 = _mid_data_in_1_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_1_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_72 = _mid_data_in_1_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_1_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_73 = _mid_data_in_1_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_1_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_74 = _mid_data_in_1_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_1_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_75 = _mid_data_in_1_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_1_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_76 = _mid_data_in_1_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_1_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_77 = _mid_data_in_1_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_1_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_78 = _mid_data_in_1_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_1_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_79 = _mid_data_in_1_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_1_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_1_tdata_T_80 = _mid_data_in_1_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_1_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_66 = _mid_data_in_1_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_1_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_67 = _mid_data_in_1_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_1_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_68 = _mid_data_in_1_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_1_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_69 = _mid_data_in_1_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_1_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_70 = _mid_data_in_1_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_1_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_71 = _mid_data_in_1_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_1_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_72 = _mid_data_in_1_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_1_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_73 = _mid_data_in_1_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_1_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_74 = _mid_data_in_1_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_1_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_75 = _mid_data_in_1_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_1_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_76 = _mid_data_in_1_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_1_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_77 = _mid_data_in_1_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_1_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_78 = _mid_data_in_1_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_1_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_79 = _mid_data_in_1_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_1_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_1_tkeep_T_80 = _mid_data_in_1_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_1_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_5 = _T_8 < 32'h10 ? _mid_data_in_1_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_6 = _T_8 < 32'h10 & _mid_data_in_1_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_1_tdata = 32'h1 >= mid_count ? _GEN_5 : mid_m_axis_tdata[63:32]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_1_tkeep = 32'h1 >= mid_count ? _GEN_6 : mid_m_axis_tkeep[1]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_12 = 32'h2 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_2_tdata_T_3 = 32'h0 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_7 = 32'h1 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_11 = 32'h2 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_15 = 32'h3 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_19 = 32'h4 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_23 = 32'h5 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_27 = 32'h6 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_31 = 32'h7 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_35 = 32'h8 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_39 = 32'h9 == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_43 = 32'ha == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_47 = 32'hb == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_51 = 32'hc == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_55 = 32'hd == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_59 = 32'he == _T_12; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_2_tdata_T_63 = 32'hf == _T_12; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_2_tdata_T_65 = _mid_data_in_2_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_66 = _mid_data_in_2_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_2_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_67 = _mid_data_in_2_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_2_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_68 = _mid_data_in_2_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_2_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_69 = _mid_data_in_2_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_2_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_70 = _mid_data_in_2_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_2_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_71 = _mid_data_in_2_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_2_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_72 = _mid_data_in_2_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_2_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_73 = _mid_data_in_2_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_2_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_74 = _mid_data_in_2_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_2_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_75 = _mid_data_in_2_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_2_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_76 = _mid_data_in_2_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_2_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_77 = _mid_data_in_2_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_2_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_78 = _mid_data_in_2_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_2_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_79 = _mid_data_in_2_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_2_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_2_tdata_T_80 = _mid_data_in_2_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_2_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_66 = _mid_data_in_2_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_2_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_67 = _mid_data_in_2_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_2_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_68 = _mid_data_in_2_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_2_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_69 = _mid_data_in_2_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_2_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_70 = _mid_data_in_2_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_2_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_71 = _mid_data_in_2_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_2_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_72 = _mid_data_in_2_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_2_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_73 = _mid_data_in_2_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_2_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_74 = _mid_data_in_2_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_2_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_75 = _mid_data_in_2_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_2_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_76 = _mid_data_in_2_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_2_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_77 = _mid_data_in_2_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_2_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_78 = _mid_data_in_2_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_2_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_79 = _mid_data_in_2_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_2_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_2_tkeep_T_80 = _mid_data_in_2_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_2_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_9 = _T_12 < 32'h10 ? _mid_data_in_2_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_10 = _T_12 < 32'h10 & _mid_data_in_2_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_2_tdata = 32'h2 >= mid_count ? _GEN_9 : mid_m_axis_tdata[95:64]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_2_tkeep = 32'h2 >= mid_count ? _GEN_10 : mid_m_axis_tkeep[2]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_16 = 32'h3 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_3_tdata_T_3 = 32'h0 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_7 = 32'h1 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_11 = 32'h2 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_15 = 32'h3 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_19 = 32'h4 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_23 = 32'h5 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_27 = 32'h6 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_31 = 32'h7 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_35 = 32'h8 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_39 = 32'h9 == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_43 = 32'ha == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_47 = 32'hb == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_51 = 32'hc == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_55 = 32'hd == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_59 = 32'he == _T_16; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_3_tdata_T_63 = 32'hf == _T_16; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_3_tdata_T_65 = _mid_data_in_3_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_66 = _mid_data_in_3_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_3_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_67 = _mid_data_in_3_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_3_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_68 = _mid_data_in_3_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_3_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_69 = _mid_data_in_3_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_3_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_70 = _mid_data_in_3_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_3_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_71 = _mid_data_in_3_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_3_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_72 = _mid_data_in_3_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_3_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_73 = _mid_data_in_3_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_3_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_74 = _mid_data_in_3_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_3_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_75 = _mid_data_in_3_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_3_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_76 = _mid_data_in_3_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_3_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_77 = _mid_data_in_3_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_3_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_78 = _mid_data_in_3_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_3_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_79 = _mid_data_in_3_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_3_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_3_tdata_T_80 = _mid_data_in_3_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_3_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_66 = _mid_data_in_3_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_3_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_67 = _mid_data_in_3_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_3_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_68 = _mid_data_in_3_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_3_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_69 = _mid_data_in_3_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_3_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_70 = _mid_data_in_3_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_3_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_71 = _mid_data_in_3_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_3_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_72 = _mid_data_in_3_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_3_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_73 = _mid_data_in_3_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_3_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_74 = _mid_data_in_3_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_3_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_75 = _mid_data_in_3_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_3_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_76 = _mid_data_in_3_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_3_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_77 = _mid_data_in_3_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_3_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_78 = _mid_data_in_3_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_3_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_79 = _mid_data_in_3_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_3_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_3_tkeep_T_80 = _mid_data_in_3_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_3_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_13 = _T_16 < 32'h10 ? _mid_data_in_3_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_14 = _T_16 < 32'h10 & _mid_data_in_3_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_3_tdata = 32'h3 >= mid_count ? _GEN_13 : mid_m_axis_tdata[127:96]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_3_tkeep = 32'h3 >= mid_count ? _GEN_14 : mid_m_axis_tkeep[3]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_20 = 32'h4 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_4_tdata_T_3 = 32'h0 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_7 = 32'h1 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_11 = 32'h2 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_15 = 32'h3 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_19 = 32'h4 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_23 = 32'h5 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_27 = 32'h6 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_31 = 32'h7 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_35 = 32'h8 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_39 = 32'h9 == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_43 = 32'ha == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_47 = 32'hb == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_51 = 32'hc == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_55 = 32'hd == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_59 = 32'he == _T_20; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_4_tdata_T_63 = 32'hf == _T_20; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_4_tdata_T_65 = _mid_data_in_4_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_66 = _mid_data_in_4_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_4_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_67 = _mid_data_in_4_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_4_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_68 = _mid_data_in_4_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_4_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_69 = _mid_data_in_4_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_4_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_70 = _mid_data_in_4_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_4_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_71 = _mid_data_in_4_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_4_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_72 = _mid_data_in_4_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_4_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_73 = _mid_data_in_4_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_4_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_74 = _mid_data_in_4_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_4_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_75 = _mid_data_in_4_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_4_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_76 = _mid_data_in_4_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_4_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_77 = _mid_data_in_4_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_4_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_78 = _mid_data_in_4_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_4_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_79 = _mid_data_in_4_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_4_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_4_tdata_T_80 = _mid_data_in_4_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_4_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_66 = _mid_data_in_4_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_4_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_67 = _mid_data_in_4_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_4_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_68 = _mid_data_in_4_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_4_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_69 = _mid_data_in_4_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_4_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_70 = _mid_data_in_4_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_4_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_71 = _mid_data_in_4_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_4_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_72 = _mid_data_in_4_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_4_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_73 = _mid_data_in_4_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_4_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_74 = _mid_data_in_4_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_4_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_75 = _mid_data_in_4_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_4_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_76 = _mid_data_in_4_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_4_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_77 = _mid_data_in_4_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_4_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_78 = _mid_data_in_4_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_4_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_79 = _mid_data_in_4_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_4_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_4_tkeep_T_80 = _mid_data_in_4_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_4_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_17 = _T_20 < 32'h10 ? _mid_data_in_4_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_18 = _T_20 < 32'h10 & _mid_data_in_4_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_4_tdata = 32'h4 >= mid_count ? _GEN_17 : mid_m_axis_tdata[159:128]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_4_tkeep = 32'h4 >= mid_count ? _GEN_18 : mid_m_axis_tkeep[4]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_24 = 32'h5 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_5_tdata_T_3 = 32'h0 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_7 = 32'h1 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_11 = 32'h2 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_15 = 32'h3 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_19 = 32'h4 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_23 = 32'h5 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_27 = 32'h6 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_31 = 32'h7 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_35 = 32'h8 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_39 = 32'h9 == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_43 = 32'ha == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_47 = 32'hb == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_51 = 32'hc == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_55 = 32'hd == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_59 = 32'he == _T_24; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_5_tdata_T_63 = 32'hf == _T_24; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_5_tdata_T_65 = _mid_data_in_5_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_66 = _mid_data_in_5_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_5_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_67 = _mid_data_in_5_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_5_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_68 = _mid_data_in_5_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_5_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_69 = _mid_data_in_5_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_5_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_70 = _mid_data_in_5_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_5_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_71 = _mid_data_in_5_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_5_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_72 = _mid_data_in_5_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_5_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_73 = _mid_data_in_5_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_5_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_74 = _mid_data_in_5_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_5_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_75 = _mid_data_in_5_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_5_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_76 = _mid_data_in_5_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_5_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_77 = _mid_data_in_5_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_5_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_78 = _mid_data_in_5_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_5_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_79 = _mid_data_in_5_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_5_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_5_tdata_T_80 = _mid_data_in_5_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_5_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_66 = _mid_data_in_5_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_5_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_67 = _mid_data_in_5_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_5_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_68 = _mid_data_in_5_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_5_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_69 = _mid_data_in_5_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_5_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_70 = _mid_data_in_5_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_5_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_71 = _mid_data_in_5_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_5_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_72 = _mid_data_in_5_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_5_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_73 = _mid_data_in_5_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_5_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_74 = _mid_data_in_5_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_5_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_75 = _mid_data_in_5_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_5_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_76 = _mid_data_in_5_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_5_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_77 = _mid_data_in_5_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_5_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_78 = _mid_data_in_5_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_5_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_79 = _mid_data_in_5_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_5_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_5_tkeep_T_80 = _mid_data_in_5_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_5_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_21 = _T_24 < 32'h10 ? _mid_data_in_5_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_22 = _T_24 < 32'h10 & _mid_data_in_5_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_5_tdata = 32'h5 >= mid_count ? _GEN_21 : mid_m_axis_tdata[191:160]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_5_tkeep = 32'h5 >= mid_count ? _GEN_22 : mid_m_axis_tkeep[5]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_28 = 32'h6 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_6_tdata_T_3 = 32'h0 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_7 = 32'h1 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_11 = 32'h2 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_15 = 32'h3 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_19 = 32'h4 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_23 = 32'h5 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_27 = 32'h6 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_31 = 32'h7 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_35 = 32'h8 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_39 = 32'h9 == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_43 = 32'ha == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_47 = 32'hb == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_51 = 32'hc == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_55 = 32'hd == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_59 = 32'he == _T_28; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_6_tdata_T_63 = 32'hf == _T_28; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_6_tdata_T_65 = _mid_data_in_6_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_66 = _mid_data_in_6_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_6_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_67 = _mid_data_in_6_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_6_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_68 = _mid_data_in_6_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_6_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_69 = _mid_data_in_6_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_6_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_70 = _mid_data_in_6_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_6_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_71 = _mid_data_in_6_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_6_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_72 = _mid_data_in_6_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_6_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_73 = _mid_data_in_6_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_6_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_74 = _mid_data_in_6_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_6_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_75 = _mid_data_in_6_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_6_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_76 = _mid_data_in_6_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_6_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_77 = _mid_data_in_6_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_6_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_78 = _mid_data_in_6_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_6_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_79 = _mid_data_in_6_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_6_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_6_tdata_T_80 = _mid_data_in_6_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_6_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_66 = _mid_data_in_6_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_6_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_67 = _mid_data_in_6_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_6_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_68 = _mid_data_in_6_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_6_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_69 = _mid_data_in_6_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_6_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_70 = _mid_data_in_6_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_6_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_71 = _mid_data_in_6_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_6_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_72 = _mid_data_in_6_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_6_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_73 = _mid_data_in_6_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_6_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_74 = _mid_data_in_6_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_6_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_75 = _mid_data_in_6_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_6_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_76 = _mid_data_in_6_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_6_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_77 = _mid_data_in_6_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_6_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_78 = _mid_data_in_6_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_6_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_79 = _mid_data_in_6_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_6_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_6_tkeep_T_80 = _mid_data_in_6_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_6_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_25 = _T_28 < 32'h10 ? _mid_data_in_6_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_26 = _T_28 < 32'h10 & _mid_data_in_6_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_6_tdata = 32'h6 >= mid_count ? _GEN_25 : mid_m_axis_tdata[223:192]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_6_tkeep = 32'h6 >= mid_count ? _GEN_26 : mid_m_axis_tkeep[6]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_32 = 32'h7 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_7_tdata_T_3 = 32'h0 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_7 = 32'h1 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_11 = 32'h2 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_15 = 32'h3 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_19 = 32'h4 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_23 = 32'h5 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_27 = 32'h6 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_31 = 32'h7 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_35 = 32'h8 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_39 = 32'h9 == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_43 = 32'ha == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_47 = 32'hb == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_51 = 32'hc == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_55 = 32'hd == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_59 = 32'he == _T_32; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_7_tdata_T_63 = 32'hf == _T_32; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_7_tdata_T_65 = _mid_data_in_7_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_66 = _mid_data_in_7_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_7_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_67 = _mid_data_in_7_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_7_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_68 = _mid_data_in_7_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_7_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_69 = _mid_data_in_7_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_7_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_70 = _mid_data_in_7_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_7_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_71 = _mid_data_in_7_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_7_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_72 = _mid_data_in_7_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_7_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_73 = _mid_data_in_7_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_7_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_74 = _mid_data_in_7_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_7_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_75 = _mid_data_in_7_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_7_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_76 = _mid_data_in_7_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_7_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_77 = _mid_data_in_7_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_7_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_78 = _mid_data_in_7_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_7_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_79 = _mid_data_in_7_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_7_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_7_tdata_T_80 = _mid_data_in_7_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_7_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_66 = _mid_data_in_7_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_7_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_67 = _mid_data_in_7_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_7_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_68 = _mid_data_in_7_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_7_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_69 = _mid_data_in_7_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_7_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_70 = _mid_data_in_7_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_7_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_71 = _mid_data_in_7_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_7_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_72 = _mid_data_in_7_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_7_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_73 = _mid_data_in_7_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_7_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_74 = _mid_data_in_7_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_7_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_75 = _mid_data_in_7_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_7_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_76 = _mid_data_in_7_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_7_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_77 = _mid_data_in_7_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_7_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_78 = _mid_data_in_7_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_7_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_79 = _mid_data_in_7_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_7_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_7_tkeep_T_80 = _mid_data_in_7_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_7_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_29 = _T_32 < 32'h10 ? _mid_data_in_7_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_30 = _T_32 < 32'h10 & _mid_data_in_7_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_7_tdata = 32'h7 >= mid_count ? _GEN_29 : mid_m_axis_tdata[255:224]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_7_tkeep = 32'h7 >= mid_count ? _GEN_30 : mid_m_axis_tkeep[7]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_36 = 32'h8 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_8_tdata_T_3 = 32'h0 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_7 = 32'h1 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_11 = 32'h2 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_15 = 32'h3 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_19 = 32'h4 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_23 = 32'h5 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_27 = 32'h6 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_31 = 32'h7 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_35 = 32'h8 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_39 = 32'h9 == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_43 = 32'ha == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_47 = 32'hb == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_51 = 32'hc == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_55 = 32'hd == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_59 = 32'he == _T_36; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_8_tdata_T_63 = 32'hf == _T_36; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_8_tdata_T_65 = _mid_data_in_8_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_66 = _mid_data_in_8_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_8_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_67 = _mid_data_in_8_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_8_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_68 = _mid_data_in_8_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_8_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_69 = _mid_data_in_8_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_8_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_70 = _mid_data_in_8_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_8_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_71 = _mid_data_in_8_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_8_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_72 = _mid_data_in_8_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_8_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_73 = _mid_data_in_8_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_8_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_74 = _mid_data_in_8_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_8_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_75 = _mid_data_in_8_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_8_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_76 = _mid_data_in_8_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_8_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_77 = _mid_data_in_8_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_8_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_78 = _mid_data_in_8_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_8_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_79 = _mid_data_in_8_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_8_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_8_tdata_T_80 = _mid_data_in_8_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_8_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_66 = _mid_data_in_8_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_8_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_67 = _mid_data_in_8_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_8_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_68 = _mid_data_in_8_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_8_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_69 = _mid_data_in_8_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_8_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_70 = _mid_data_in_8_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_8_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_71 = _mid_data_in_8_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_8_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_72 = _mid_data_in_8_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_8_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_73 = _mid_data_in_8_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_8_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_74 = _mid_data_in_8_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_8_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_75 = _mid_data_in_8_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_8_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_76 = _mid_data_in_8_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_8_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_77 = _mid_data_in_8_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_8_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_78 = _mid_data_in_8_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_8_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_79 = _mid_data_in_8_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_8_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_8_tkeep_T_80 = _mid_data_in_8_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_8_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_33 = _T_36 < 32'h10 ? _mid_data_in_8_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_34 = _T_36 < 32'h10 & _mid_data_in_8_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_8_tdata = 32'h8 >= mid_count ? _GEN_33 : mid_m_axis_tdata[287:256]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_8_tkeep = 32'h8 >= mid_count ? _GEN_34 : mid_m_axis_tkeep[8]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_40 = 32'h9 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_9_tdata_T_3 = 32'h0 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_7 = 32'h1 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_11 = 32'h2 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_15 = 32'h3 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_19 = 32'h4 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_23 = 32'h5 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_27 = 32'h6 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_31 = 32'h7 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_35 = 32'h8 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_39 = 32'h9 == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_43 = 32'ha == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_47 = 32'hb == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_51 = 32'hc == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_55 = 32'hd == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_59 = 32'he == _T_40; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_9_tdata_T_63 = 32'hf == _T_40; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_9_tdata_T_65 = _mid_data_in_9_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_66 = _mid_data_in_9_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_9_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_67 = _mid_data_in_9_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_9_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_68 = _mid_data_in_9_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_9_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_69 = _mid_data_in_9_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_9_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_70 = _mid_data_in_9_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_9_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_71 = _mid_data_in_9_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_9_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_72 = _mid_data_in_9_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_9_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_73 = _mid_data_in_9_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_9_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_74 = _mid_data_in_9_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_9_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_75 = _mid_data_in_9_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_9_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_76 = _mid_data_in_9_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_9_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_77 = _mid_data_in_9_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_9_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_78 = _mid_data_in_9_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_9_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_79 = _mid_data_in_9_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_9_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_9_tdata_T_80 = _mid_data_in_9_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_9_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_66 = _mid_data_in_9_tdata_T_59 ? sorted_in_m_axis_tkeep[14] : _mid_data_in_9_tdata_T_63
     & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_67 = _mid_data_in_9_tdata_T_55 ? sorted_in_m_axis_tkeep[13] : _mid_data_in_9_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_68 = _mid_data_in_9_tdata_T_51 ? sorted_in_m_axis_tkeep[12] : _mid_data_in_9_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_69 = _mid_data_in_9_tdata_T_47 ? sorted_in_m_axis_tkeep[11] : _mid_data_in_9_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_70 = _mid_data_in_9_tdata_T_43 ? sorted_in_m_axis_tkeep[10] : _mid_data_in_9_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_71 = _mid_data_in_9_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_9_tkeep_T_70; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_72 = _mid_data_in_9_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_9_tkeep_T_71; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_73 = _mid_data_in_9_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_9_tkeep_T_72; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_74 = _mid_data_in_9_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_9_tkeep_T_73; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_75 = _mid_data_in_9_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_9_tkeep_T_74; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_76 = _mid_data_in_9_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_9_tkeep_T_75; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_77 = _mid_data_in_9_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_9_tkeep_T_76; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_78 = _mid_data_in_9_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_9_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_79 = _mid_data_in_9_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_9_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_9_tkeep_T_80 = _mid_data_in_9_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_9_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_37 = _T_40 < 32'h10 ? _mid_data_in_9_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_38 = _T_40 < 32'h10 & _mid_data_in_9_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_9_tdata = 32'h9 >= mid_count ? _GEN_37 : mid_m_axis_tdata[319:288]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_9_tkeep = 32'h9 >= mid_count ? _GEN_38 : mid_m_axis_tkeep[9]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_44 = 32'ha - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_10_tdata_T_3 = 32'h0 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_7 = 32'h1 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_11 = 32'h2 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_15 = 32'h3 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_19 = 32'h4 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_23 = 32'h5 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_27 = 32'h6 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_31 = 32'h7 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_35 = 32'h8 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_39 = 32'h9 == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_43 = 32'ha == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_47 = 32'hb == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_51 = 32'hc == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_55 = 32'hd == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_59 = 32'he == _T_44; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_10_tdata_T_63 = 32'hf == _T_44; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_10_tdata_T_65 = _mid_data_in_10_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_66 = _mid_data_in_10_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_10_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_67 = _mid_data_in_10_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_10_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_68 = _mid_data_in_10_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_10_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_69 = _mid_data_in_10_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_10_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_70 = _mid_data_in_10_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_10_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_71 = _mid_data_in_10_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_10_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_72 = _mid_data_in_10_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_10_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_73 = _mid_data_in_10_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_10_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_74 = _mid_data_in_10_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_10_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_75 = _mid_data_in_10_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_10_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_76 = _mid_data_in_10_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_10_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_77 = _mid_data_in_10_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_10_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_78 = _mid_data_in_10_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_10_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_79 = _mid_data_in_10_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_10_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_10_tdata_T_80 = _mid_data_in_10_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_10_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_66 = _mid_data_in_10_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_10_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_67 = _mid_data_in_10_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_10_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_68 = _mid_data_in_10_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_10_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_69 = _mid_data_in_10_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_10_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_70 = _mid_data_in_10_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_10_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_71 = _mid_data_in_10_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_10_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_72 = _mid_data_in_10_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_10_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_73 = _mid_data_in_10_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_10_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_74 = _mid_data_in_10_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_10_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_75 = _mid_data_in_10_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_10_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_76 = _mid_data_in_10_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_10_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_77 = _mid_data_in_10_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_10_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_78 = _mid_data_in_10_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_10_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_79 = _mid_data_in_10_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_10_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_10_tkeep_T_80 = _mid_data_in_10_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_10_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_41 = _T_44 < 32'h10 ? _mid_data_in_10_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_42 = _T_44 < 32'h10 & _mid_data_in_10_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_10_tdata = 32'ha >= mid_count ? _GEN_41 : mid_m_axis_tdata[351:320]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_10_tkeep = 32'ha >= mid_count ? _GEN_42 : mid_m_axis_tkeep[10]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_48 = 32'hb - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_11_tdata_T_3 = 32'h0 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_7 = 32'h1 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_11 = 32'h2 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_15 = 32'h3 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_19 = 32'h4 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_23 = 32'h5 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_27 = 32'h6 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_31 = 32'h7 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_35 = 32'h8 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_39 = 32'h9 == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_43 = 32'ha == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_47 = 32'hb == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_51 = 32'hc == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_55 = 32'hd == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_59 = 32'he == _T_48; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_11_tdata_T_63 = 32'hf == _T_48; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_11_tdata_T_65 = _mid_data_in_11_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_66 = _mid_data_in_11_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_11_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_67 = _mid_data_in_11_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_11_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_68 = _mid_data_in_11_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_11_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_69 = _mid_data_in_11_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_11_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_70 = _mid_data_in_11_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_11_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_71 = _mid_data_in_11_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_11_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_72 = _mid_data_in_11_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_11_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_73 = _mid_data_in_11_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_11_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_74 = _mid_data_in_11_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_11_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_75 = _mid_data_in_11_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_11_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_76 = _mid_data_in_11_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_11_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_77 = _mid_data_in_11_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_11_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_78 = _mid_data_in_11_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_11_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_79 = _mid_data_in_11_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_11_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_11_tdata_T_80 = _mid_data_in_11_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_11_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_66 = _mid_data_in_11_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_11_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_67 = _mid_data_in_11_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_11_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_68 = _mid_data_in_11_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_11_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_69 = _mid_data_in_11_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_11_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_70 = _mid_data_in_11_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_11_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_71 = _mid_data_in_11_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_11_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_72 = _mid_data_in_11_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_11_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_73 = _mid_data_in_11_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_11_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_74 = _mid_data_in_11_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_11_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_75 = _mid_data_in_11_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_11_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_76 = _mid_data_in_11_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_11_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_77 = _mid_data_in_11_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_11_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_78 = _mid_data_in_11_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_11_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_79 = _mid_data_in_11_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_11_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_11_tkeep_T_80 = _mid_data_in_11_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_11_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_45 = _T_48 < 32'h10 ? _mid_data_in_11_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_46 = _T_48 < 32'h10 & _mid_data_in_11_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_11_tdata = 32'hb >= mid_count ? _GEN_45 : mid_m_axis_tdata[383:352]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_11_tkeep = 32'hb >= mid_count ? _GEN_46 : mid_m_axis_tkeep[11]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_52 = 32'hc - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_12_tdata_T_3 = 32'h0 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_7 = 32'h1 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_11 = 32'h2 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_15 = 32'h3 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_19 = 32'h4 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_23 = 32'h5 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_27 = 32'h6 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_31 = 32'h7 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_35 = 32'h8 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_39 = 32'h9 == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_43 = 32'ha == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_47 = 32'hb == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_51 = 32'hc == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_55 = 32'hd == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_59 = 32'he == _T_52; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_12_tdata_T_63 = 32'hf == _T_52; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_12_tdata_T_65 = _mid_data_in_12_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_66 = _mid_data_in_12_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_12_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_67 = _mid_data_in_12_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_12_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_68 = _mid_data_in_12_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_12_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_69 = _mid_data_in_12_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_12_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_70 = _mid_data_in_12_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_12_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_71 = _mid_data_in_12_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_12_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_72 = _mid_data_in_12_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_12_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_73 = _mid_data_in_12_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_12_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_74 = _mid_data_in_12_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_12_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_75 = _mid_data_in_12_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_12_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_76 = _mid_data_in_12_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_12_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_77 = _mid_data_in_12_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_12_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_78 = _mid_data_in_12_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_12_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_79 = _mid_data_in_12_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_12_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_12_tdata_T_80 = _mid_data_in_12_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_12_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_66 = _mid_data_in_12_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_12_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_67 = _mid_data_in_12_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_12_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_68 = _mid_data_in_12_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_12_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_69 = _mid_data_in_12_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_12_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_70 = _mid_data_in_12_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_12_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_71 = _mid_data_in_12_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_12_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_72 = _mid_data_in_12_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_12_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_73 = _mid_data_in_12_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_12_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_74 = _mid_data_in_12_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_12_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_75 = _mid_data_in_12_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_12_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_76 = _mid_data_in_12_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_12_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_77 = _mid_data_in_12_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_12_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_78 = _mid_data_in_12_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_12_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_79 = _mid_data_in_12_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_12_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_12_tkeep_T_80 = _mid_data_in_12_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_12_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_49 = _T_52 < 32'h10 ? _mid_data_in_12_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_50 = _T_52 < 32'h10 & _mid_data_in_12_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_12_tdata = 32'hc >= mid_count ? _GEN_49 : mid_m_axis_tdata[415:384]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_12_tkeep = 32'hc >= mid_count ? _GEN_50 : mid_m_axis_tkeep[12]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_56 = 32'hd - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_13_tdata_T_3 = 32'h0 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_7 = 32'h1 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_11 = 32'h2 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_15 = 32'h3 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_19 = 32'h4 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_23 = 32'h5 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_27 = 32'h6 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_31 = 32'h7 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_35 = 32'h8 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_39 = 32'h9 == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_43 = 32'ha == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_47 = 32'hb == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_51 = 32'hc == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_55 = 32'hd == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_59 = 32'he == _T_56; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_13_tdata_T_63 = 32'hf == _T_56; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_13_tdata_T_65 = _mid_data_in_13_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_66 = _mid_data_in_13_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_13_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_67 = _mid_data_in_13_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_13_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_68 = _mid_data_in_13_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_13_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_69 = _mid_data_in_13_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_13_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_70 = _mid_data_in_13_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_13_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_71 = _mid_data_in_13_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_13_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_72 = _mid_data_in_13_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_13_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_73 = _mid_data_in_13_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_13_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_74 = _mid_data_in_13_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_13_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_75 = _mid_data_in_13_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_13_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_76 = _mid_data_in_13_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_13_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_77 = _mid_data_in_13_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_13_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_78 = _mid_data_in_13_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_13_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_79 = _mid_data_in_13_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_13_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_13_tdata_T_80 = _mid_data_in_13_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_13_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_66 = _mid_data_in_13_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_13_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_67 = _mid_data_in_13_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_13_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_68 = _mid_data_in_13_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_13_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_69 = _mid_data_in_13_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_13_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_70 = _mid_data_in_13_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_13_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_71 = _mid_data_in_13_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_13_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_72 = _mid_data_in_13_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_13_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_73 = _mid_data_in_13_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_13_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_74 = _mid_data_in_13_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_13_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_75 = _mid_data_in_13_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_13_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_76 = _mid_data_in_13_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_13_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_77 = _mid_data_in_13_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_13_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_78 = _mid_data_in_13_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_13_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_79 = _mid_data_in_13_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_13_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_13_tkeep_T_80 = _mid_data_in_13_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_13_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_53 = _T_56 < 32'h10 ? _mid_data_in_13_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_54 = _T_56 < 32'h10 & _mid_data_in_13_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_13_tdata = 32'hd >= mid_count ? _GEN_53 : mid_m_axis_tdata[447:416]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_13_tkeep = 32'hd >= mid_count ? _GEN_54 : mid_m_axis_tkeep[13]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_60 = 32'he - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_14_tdata_T_3 = 32'h0 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_7 = 32'h1 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_11 = 32'h2 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_15 = 32'h3 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_19 = 32'h4 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_23 = 32'h5 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_27 = 32'h6 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_31 = 32'h7 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_35 = 32'h8 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_39 = 32'h9 == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_43 = 32'ha == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_47 = 32'hb == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_51 = 32'hc == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_55 = 32'hd == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_59 = 32'he == _T_60; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_14_tdata_T_63 = 32'hf == _T_60; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_14_tdata_T_65 = _mid_data_in_14_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_66 = _mid_data_in_14_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_14_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_67 = _mid_data_in_14_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_14_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_68 = _mid_data_in_14_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_14_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_69 = _mid_data_in_14_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_14_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_70 = _mid_data_in_14_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_14_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_71 = _mid_data_in_14_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_14_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_72 = _mid_data_in_14_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_14_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_73 = _mid_data_in_14_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_14_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_74 = _mid_data_in_14_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_14_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_75 = _mid_data_in_14_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_14_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_76 = _mid_data_in_14_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_14_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_77 = _mid_data_in_14_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_14_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_78 = _mid_data_in_14_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_14_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_79 = _mid_data_in_14_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_14_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_14_tdata_T_80 = _mid_data_in_14_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_14_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_66 = _mid_data_in_14_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_14_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_67 = _mid_data_in_14_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_14_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_68 = _mid_data_in_14_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_14_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_69 = _mid_data_in_14_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_14_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_70 = _mid_data_in_14_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_14_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_71 = _mid_data_in_14_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_14_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_72 = _mid_data_in_14_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_14_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_73 = _mid_data_in_14_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_14_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_74 = _mid_data_in_14_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_14_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_75 = _mid_data_in_14_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_14_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_76 = _mid_data_in_14_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_14_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_77 = _mid_data_in_14_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_14_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_78 = _mid_data_in_14_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_14_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_79 = _mid_data_in_14_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_14_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_14_tkeep_T_80 = _mid_data_in_14_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_14_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_57 = _T_60 < 32'h10 ? _mid_data_in_14_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_58 = _T_60 < 32'h10 & _mid_data_in_14_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_14_tdata = 32'he >= mid_count ? _GEN_57 : mid_m_axis_tdata[479:448]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_14_tkeep = 32'he >= mid_count ? _GEN_58 : mid_m_axis_tkeep[14]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_64 = 32'hf - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_15_tdata_T_3 = 32'h0 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_7 = 32'h1 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_11 = 32'h2 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_15 = 32'h3 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_19 = 32'h4 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_23 = 32'h5 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_27 = 32'h6 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_31 = 32'h7 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_35 = 32'h8 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_39 = 32'h9 == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_43 = 32'ha == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_47 = 32'hb == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_51 = 32'hc == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_55 = 32'hd == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_59 = 32'he == _T_64; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_15_tdata_T_63 = 32'hf == _T_64; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_15_tdata_T_65 = _mid_data_in_15_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_66 = _mid_data_in_15_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_15_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_67 = _mid_data_in_15_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_15_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_68 = _mid_data_in_15_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_15_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_69 = _mid_data_in_15_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_15_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_70 = _mid_data_in_15_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_15_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_71 = _mid_data_in_15_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_15_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_72 = _mid_data_in_15_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_15_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_73 = _mid_data_in_15_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_15_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_74 = _mid_data_in_15_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_15_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_75 = _mid_data_in_15_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_15_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_76 = _mid_data_in_15_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_15_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_77 = _mid_data_in_15_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_15_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_78 = _mid_data_in_15_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_15_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_79 = _mid_data_in_15_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_15_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_15_tdata_T_80 = _mid_data_in_15_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_15_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_66 = _mid_data_in_15_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_15_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_67 = _mid_data_in_15_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_15_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_68 = _mid_data_in_15_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_15_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_69 = _mid_data_in_15_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_15_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_70 = _mid_data_in_15_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_15_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_71 = _mid_data_in_15_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_15_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_72 = _mid_data_in_15_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_15_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_73 = _mid_data_in_15_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_15_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_74 = _mid_data_in_15_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_15_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_75 = _mid_data_in_15_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_15_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_76 = _mid_data_in_15_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_15_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_77 = _mid_data_in_15_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_15_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_78 = _mid_data_in_15_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_15_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_79 = _mid_data_in_15_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_15_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_15_tkeep_T_80 = _mid_data_in_15_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_15_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_61 = _T_64 < 32'h10 ? _mid_data_in_15_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_62 = _T_64 < 32'h10 & _mid_data_in_15_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_15_tdata = 32'hf >= mid_count ? _GEN_61 : mid_m_axis_tdata[511:480]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_15_tkeep = 32'hf >= mid_count ? _GEN_62 : mid_m_axis_tkeep[15]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_68 = 32'h10 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_16_tdata_T_3 = 32'h0 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_7 = 32'h1 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_11 = 32'h2 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_15 = 32'h3 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_19 = 32'h4 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_23 = 32'h5 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_27 = 32'h6 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_31 = 32'h7 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_35 = 32'h8 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_39 = 32'h9 == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_43 = 32'ha == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_47 = 32'hb == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_51 = 32'hc == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_55 = 32'hd == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_59 = 32'he == _T_68; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_16_tdata_T_63 = 32'hf == _T_68; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_16_tdata_T_65 = _mid_data_in_16_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_66 = _mid_data_in_16_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_16_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_67 = _mid_data_in_16_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_16_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_68 = _mid_data_in_16_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_16_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_69 = _mid_data_in_16_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_16_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_70 = _mid_data_in_16_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_16_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_71 = _mid_data_in_16_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_16_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_72 = _mid_data_in_16_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_16_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_73 = _mid_data_in_16_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_16_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_74 = _mid_data_in_16_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_16_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_75 = _mid_data_in_16_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_16_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_76 = _mid_data_in_16_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_16_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_77 = _mid_data_in_16_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_16_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_78 = _mid_data_in_16_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_16_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_79 = _mid_data_in_16_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_16_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_16_tdata_T_80 = _mid_data_in_16_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_16_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_66 = _mid_data_in_16_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_16_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_67 = _mid_data_in_16_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_16_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_68 = _mid_data_in_16_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_16_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_69 = _mid_data_in_16_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_16_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_70 = _mid_data_in_16_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_16_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_71 = _mid_data_in_16_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_16_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_72 = _mid_data_in_16_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_16_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_73 = _mid_data_in_16_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_16_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_74 = _mid_data_in_16_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_16_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_75 = _mid_data_in_16_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_16_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_76 = _mid_data_in_16_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_16_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_77 = _mid_data_in_16_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_16_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_78 = _mid_data_in_16_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_16_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_79 = _mid_data_in_16_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_16_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_16_tkeep_T_80 = _mid_data_in_16_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_16_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_65 = _T_68 < 32'h10 ? _mid_data_in_16_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_66 = _T_68 < 32'h10 & _mid_data_in_16_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_16_tdata = 32'h10 >= mid_count ? _GEN_65 : mid_m_axis_tdata[543:512]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_16_tkeep = 32'h10 >= mid_count ? _GEN_66 : mid_m_axis_tkeep[16]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_72 = 32'h11 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_17_tdata_T_3 = 32'h0 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_7 = 32'h1 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_11 = 32'h2 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_15 = 32'h3 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_19 = 32'h4 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_23 = 32'h5 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_27 = 32'h6 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_31 = 32'h7 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_35 = 32'h8 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_39 = 32'h9 == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_43 = 32'ha == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_47 = 32'hb == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_51 = 32'hc == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_55 = 32'hd == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_59 = 32'he == _T_72; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_17_tdata_T_63 = 32'hf == _T_72; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_17_tdata_T_65 = _mid_data_in_17_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_66 = _mid_data_in_17_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_17_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_67 = _mid_data_in_17_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_17_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_68 = _mid_data_in_17_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_17_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_69 = _mid_data_in_17_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_17_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_70 = _mid_data_in_17_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_17_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_71 = _mid_data_in_17_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_17_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_72 = _mid_data_in_17_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_17_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_73 = _mid_data_in_17_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_17_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_74 = _mid_data_in_17_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_17_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_75 = _mid_data_in_17_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_17_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_76 = _mid_data_in_17_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_17_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_77 = _mid_data_in_17_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_17_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_78 = _mid_data_in_17_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_17_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_79 = _mid_data_in_17_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_17_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_17_tdata_T_80 = _mid_data_in_17_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_17_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_66 = _mid_data_in_17_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_17_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_67 = _mid_data_in_17_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_17_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_68 = _mid_data_in_17_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_17_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_69 = _mid_data_in_17_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_17_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_70 = _mid_data_in_17_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_17_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_71 = _mid_data_in_17_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_17_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_72 = _mid_data_in_17_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_17_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_73 = _mid_data_in_17_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_17_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_74 = _mid_data_in_17_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_17_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_75 = _mid_data_in_17_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_17_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_76 = _mid_data_in_17_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_17_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_77 = _mid_data_in_17_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_17_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_78 = _mid_data_in_17_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_17_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_79 = _mid_data_in_17_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_17_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_17_tkeep_T_80 = _mid_data_in_17_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_17_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_69 = _T_72 < 32'h10 ? _mid_data_in_17_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_70 = _T_72 < 32'h10 & _mid_data_in_17_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_17_tdata = 32'h11 >= mid_count ? _GEN_69 : mid_m_axis_tdata[575:544]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_17_tkeep = 32'h11 >= mid_count ? _GEN_70 : mid_m_axis_tkeep[17]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_76 = 32'h12 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_18_tdata_T_3 = 32'h0 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_7 = 32'h1 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_11 = 32'h2 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_15 = 32'h3 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_19 = 32'h4 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_23 = 32'h5 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_27 = 32'h6 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_31 = 32'h7 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_35 = 32'h8 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_39 = 32'h9 == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_43 = 32'ha == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_47 = 32'hb == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_51 = 32'hc == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_55 = 32'hd == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_59 = 32'he == _T_76; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_18_tdata_T_63 = 32'hf == _T_76; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_18_tdata_T_65 = _mid_data_in_18_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_66 = _mid_data_in_18_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_18_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_67 = _mid_data_in_18_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_18_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_68 = _mid_data_in_18_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_18_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_69 = _mid_data_in_18_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_18_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_70 = _mid_data_in_18_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_18_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_71 = _mid_data_in_18_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_18_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_72 = _mid_data_in_18_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_18_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_73 = _mid_data_in_18_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_18_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_74 = _mid_data_in_18_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_18_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_75 = _mid_data_in_18_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_18_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_76 = _mid_data_in_18_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_18_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_77 = _mid_data_in_18_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_18_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_78 = _mid_data_in_18_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_18_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_79 = _mid_data_in_18_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_18_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_18_tdata_T_80 = _mid_data_in_18_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_18_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_66 = _mid_data_in_18_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_18_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_67 = _mid_data_in_18_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_18_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_68 = _mid_data_in_18_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_18_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_69 = _mid_data_in_18_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_18_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_70 = _mid_data_in_18_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_18_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_71 = _mid_data_in_18_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_18_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_72 = _mid_data_in_18_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_18_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_73 = _mid_data_in_18_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_18_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_74 = _mid_data_in_18_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_18_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_75 = _mid_data_in_18_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_18_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_76 = _mid_data_in_18_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_18_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_77 = _mid_data_in_18_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_18_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_78 = _mid_data_in_18_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_18_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_79 = _mid_data_in_18_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_18_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_18_tkeep_T_80 = _mid_data_in_18_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_18_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_73 = _T_76 < 32'h10 ? _mid_data_in_18_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_74 = _T_76 < 32'h10 & _mid_data_in_18_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_18_tdata = 32'h12 >= mid_count ? _GEN_73 : mid_m_axis_tdata[607:576]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_18_tkeep = 32'h12 >= mid_count ? _GEN_74 : mid_m_axis_tkeep[18]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_80 = 32'h13 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_19_tdata_T_3 = 32'h0 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_7 = 32'h1 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_11 = 32'h2 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_15 = 32'h3 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_19 = 32'h4 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_23 = 32'h5 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_27 = 32'h6 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_31 = 32'h7 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_35 = 32'h8 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_39 = 32'h9 == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_43 = 32'ha == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_47 = 32'hb == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_51 = 32'hc == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_55 = 32'hd == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_59 = 32'he == _T_80; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_19_tdata_T_63 = 32'hf == _T_80; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_19_tdata_T_65 = _mid_data_in_19_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_66 = _mid_data_in_19_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_19_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_67 = _mid_data_in_19_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_19_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_68 = _mid_data_in_19_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_19_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_69 = _mid_data_in_19_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_19_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_70 = _mid_data_in_19_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_19_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_71 = _mid_data_in_19_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_19_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_72 = _mid_data_in_19_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_19_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_73 = _mid_data_in_19_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_19_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_74 = _mid_data_in_19_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_19_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_75 = _mid_data_in_19_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_19_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_76 = _mid_data_in_19_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_19_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_77 = _mid_data_in_19_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_19_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_78 = _mid_data_in_19_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_19_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_79 = _mid_data_in_19_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_19_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_19_tdata_T_80 = _mid_data_in_19_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_19_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_66 = _mid_data_in_19_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_19_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_67 = _mid_data_in_19_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_19_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_68 = _mid_data_in_19_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_19_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_69 = _mid_data_in_19_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_19_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_70 = _mid_data_in_19_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_19_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_71 = _mid_data_in_19_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_19_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_72 = _mid_data_in_19_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_19_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_73 = _mid_data_in_19_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_19_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_74 = _mid_data_in_19_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_19_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_75 = _mid_data_in_19_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_19_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_76 = _mid_data_in_19_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_19_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_77 = _mid_data_in_19_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_19_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_78 = _mid_data_in_19_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_19_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_79 = _mid_data_in_19_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_19_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_19_tkeep_T_80 = _mid_data_in_19_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_19_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_77 = _T_80 < 32'h10 ? _mid_data_in_19_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_78 = _T_80 < 32'h10 & _mid_data_in_19_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_19_tdata = 32'h13 >= mid_count ? _GEN_77 : mid_m_axis_tdata[639:608]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_19_tkeep = 32'h13 >= mid_count ? _GEN_78 : mid_m_axis_tkeep[19]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_84 = 32'h14 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_20_tdata_T_3 = 32'h0 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_7 = 32'h1 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_11 = 32'h2 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_15 = 32'h3 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_19 = 32'h4 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_23 = 32'h5 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_27 = 32'h6 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_31 = 32'h7 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_35 = 32'h8 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_39 = 32'h9 == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_43 = 32'ha == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_47 = 32'hb == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_51 = 32'hc == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_55 = 32'hd == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_59 = 32'he == _T_84; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_20_tdata_T_63 = 32'hf == _T_84; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_20_tdata_T_65 = _mid_data_in_20_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_66 = _mid_data_in_20_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_20_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_67 = _mid_data_in_20_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_20_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_68 = _mid_data_in_20_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_20_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_69 = _mid_data_in_20_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_20_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_70 = _mid_data_in_20_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_20_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_71 = _mid_data_in_20_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_20_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_72 = _mid_data_in_20_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_20_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_73 = _mid_data_in_20_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_20_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_74 = _mid_data_in_20_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_20_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_75 = _mid_data_in_20_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_20_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_76 = _mid_data_in_20_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_20_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_77 = _mid_data_in_20_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_20_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_78 = _mid_data_in_20_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_20_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_79 = _mid_data_in_20_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_20_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_20_tdata_T_80 = _mid_data_in_20_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_20_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_66 = _mid_data_in_20_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_20_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_67 = _mid_data_in_20_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_20_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_68 = _mid_data_in_20_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_20_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_69 = _mid_data_in_20_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_20_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_70 = _mid_data_in_20_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_20_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_71 = _mid_data_in_20_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_20_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_72 = _mid_data_in_20_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_20_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_73 = _mid_data_in_20_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_20_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_74 = _mid_data_in_20_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_20_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_75 = _mid_data_in_20_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_20_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_76 = _mid_data_in_20_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_20_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_77 = _mid_data_in_20_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_20_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_78 = _mid_data_in_20_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_20_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_79 = _mid_data_in_20_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_20_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_20_tkeep_T_80 = _mid_data_in_20_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_20_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_81 = _T_84 < 32'h10 ? _mid_data_in_20_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_82 = _T_84 < 32'h10 & _mid_data_in_20_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_20_tdata = 32'h14 >= mid_count ? _GEN_81 : mid_m_axis_tdata[671:640]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_20_tkeep = 32'h14 >= mid_count ? _GEN_82 : mid_m_axis_tkeep[20]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_88 = 32'h15 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_21_tdata_T_3 = 32'h0 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_7 = 32'h1 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_11 = 32'h2 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_15 = 32'h3 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_19 = 32'h4 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_23 = 32'h5 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_27 = 32'h6 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_31 = 32'h7 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_35 = 32'h8 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_39 = 32'h9 == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_43 = 32'ha == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_47 = 32'hb == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_51 = 32'hc == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_55 = 32'hd == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_59 = 32'he == _T_88; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_21_tdata_T_63 = 32'hf == _T_88; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_21_tdata_T_65 = _mid_data_in_21_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_66 = _mid_data_in_21_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_21_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_67 = _mid_data_in_21_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_21_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_68 = _mid_data_in_21_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_21_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_69 = _mid_data_in_21_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_21_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_70 = _mid_data_in_21_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_21_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_71 = _mid_data_in_21_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_21_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_72 = _mid_data_in_21_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_21_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_73 = _mid_data_in_21_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_21_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_74 = _mid_data_in_21_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_21_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_75 = _mid_data_in_21_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_21_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_76 = _mid_data_in_21_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_21_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_77 = _mid_data_in_21_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_21_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_78 = _mid_data_in_21_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_21_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_79 = _mid_data_in_21_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_21_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_21_tdata_T_80 = _mid_data_in_21_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_21_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_66 = _mid_data_in_21_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_21_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_67 = _mid_data_in_21_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_21_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_68 = _mid_data_in_21_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_21_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_69 = _mid_data_in_21_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_21_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_70 = _mid_data_in_21_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_21_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_71 = _mid_data_in_21_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_21_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_72 = _mid_data_in_21_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_21_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_73 = _mid_data_in_21_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_21_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_74 = _mid_data_in_21_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_21_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_75 = _mid_data_in_21_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_21_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_76 = _mid_data_in_21_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_21_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_77 = _mid_data_in_21_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_21_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_78 = _mid_data_in_21_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_21_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_79 = _mid_data_in_21_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_21_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_21_tkeep_T_80 = _mid_data_in_21_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_21_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_85 = _T_88 < 32'h10 ? _mid_data_in_21_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_86 = _T_88 < 32'h10 & _mid_data_in_21_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_21_tdata = 32'h15 >= mid_count ? _GEN_85 : mid_m_axis_tdata[703:672]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_21_tkeep = 32'h15 >= mid_count ? _GEN_86 : mid_m_axis_tkeep[21]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_92 = 32'h16 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_22_tdata_T_3 = 32'h0 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_7 = 32'h1 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_11 = 32'h2 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_15 = 32'h3 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_19 = 32'h4 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_23 = 32'h5 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_27 = 32'h6 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_31 = 32'h7 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_35 = 32'h8 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_39 = 32'h9 == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_43 = 32'ha == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_47 = 32'hb == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_51 = 32'hc == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_55 = 32'hd == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_59 = 32'he == _T_92; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_22_tdata_T_63 = 32'hf == _T_92; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_22_tdata_T_65 = _mid_data_in_22_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_66 = _mid_data_in_22_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_22_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_67 = _mid_data_in_22_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_22_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_68 = _mid_data_in_22_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_22_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_69 = _mid_data_in_22_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_22_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_70 = _mid_data_in_22_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_22_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_71 = _mid_data_in_22_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_22_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_72 = _mid_data_in_22_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_22_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_73 = _mid_data_in_22_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_22_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_74 = _mid_data_in_22_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_22_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_75 = _mid_data_in_22_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_22_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_76 = _mid_data_in_22_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_22_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_77 = _mid_data_in_22_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_22_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_78 = _mid_data_in_22_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_22_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_79 = _mid_data_in_22_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_22_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_22_tdata_T_80 = _mid_data_in_22_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_22_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_66 = _mid_data_in_22_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_22_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_67 = _mid_data_in_22_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_22_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_68 = _mid_data_in_22_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_22_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_69 = _mid_data_in_22_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_22_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_70 = _mid_data_in_22_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_22_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_71 = _mid_data_in_22_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_22_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_72 = _mid_data_in_22_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_22_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_73 = _mid_data_in_22_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_22_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_74 = _mid_data_in_22_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_22_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_75 = _mid_data_in_22_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_22_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_76 = _mid_data_in_22_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_22_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_77 = _mid_data_in_22_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_22_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_78 = _mid_data_in_22_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_22_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_79 = _mid_data_in_22_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_22_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_22_tkeep_T_80 = _mid_data_in_22_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_22_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_89 = _T_92 < 32'h10 ? _mid_data_in_22_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_90 = _T_92 < 32'h10 & _mid_data_in_22_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_22_tdata = 32'h16 >= mid_count ? _GEN_89 : mid_m_axis_tdata[735:704]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_22_tkeep = 32'h16 >= mid_count ? _GEN_90 : mid_m_axis_tkeep[22]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_96 = 32'h17 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_23_tdata_T_3 = 32'h0 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_7 = 32'h1 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_11 = 32'h2 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_15 = 32'h3 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_19 = 32'h4 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_23 = 32'h5 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_27 = 32'h6 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_31 = 32'h7 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_35 = 32'h8 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_39 = 32'h9 == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_43 = 32'ha == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_47 = 32'hb == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_51 = 32'hc == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_55 = 32'hd == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_59 = 32'he == _T_96; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_23_tdata_T_63 = 32'hf == _T_96; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_23_tdata_T_65 = _mid_data_in_23_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_66 = _mid_data_in_23_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_23_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_67 = _mid_data_in_23_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_23_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_68 = _mid_data_in_23_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_23_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_69 = _mid_data_in_23_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_23_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_70 = _mid_data_in_23_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_23_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_71 = _mid_data_in_23_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_23_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_72 = _mid_data_in_23_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_23_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_73 = _mid_data_in_23_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_23_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_74 = _mid_data_in_23_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_23_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_75 = _mid_data_in_23_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_23_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_76 = _mid_data_in_23_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_23_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_77 = _mid_data_in_23_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_23_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_78 = _mid_data_in_23_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_23_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_79 = _mid_data_in_23_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_23_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_23_tdata_T_80 = _mid_data_in_23_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_23_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_66 = _mid_data_in_23_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_23_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_67 = _mid_data_in_23_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_23_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_68 = _mid_data_in_23_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_23_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_69 = _mid_data_in_23_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_23_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_70 = _mid_data_in_23_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_23_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_71 = _mid_data_in_23_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_23_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_72 = _mid_data_in_23_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_23_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_73 = _mid_data_in_23_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_23_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_74 = _mid_data_in_23_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_23_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_75 = _mid_data_in_23_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_23_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_76 = _mid_data_in_23_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_23_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_77 = _mid_data_in_23_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_23_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_78 = _mid_data_in_23_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_23_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_79 = _mid_data_in_23_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_23_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_23_tkeep_T_80 = _mid_data_in_23_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_23_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_93 = _T_96 < 32'h10 ? _mid_data_in_23_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_94 = _T_96 < 32'h10 & _mid_data_in_23_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_23_tdata = 32'h17 >= mid_count ? _GEN_93 : mid_m_axis_tdata[767:736]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_23_tkeep = 32'h17 >= mid_count ? _GEN_94 : mid_m_axis_tkeep[23]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_100 = 32'h18 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_24_tdata_T_3 = 32'h0 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_7 = 32'h1 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_11 = 32'h2 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_15 = 32'h3 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_19 = 32'h4 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_23 = 32'h5 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_27 = 32'h6 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_31 = 32'h7 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_35 = 32'h8 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_39 = 32'h9 == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_43 = 32'ha == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_47 = 32'hb == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_51 = 32'hc == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_55 = 32'hd == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_59 = 32'he == _T_100; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_24_tdata_T_63 = 32'hf == _T_100; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_24_tdata_T_65 = _mid_data_in_24_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_66 = _mid_data_in_24_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_24_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_67 = _mid_data_in_24_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_24_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_68 = _mid_data_in_24_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_24_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_69 = _mid_data_in_24_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_24_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_70 = _mid_data_in_24_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_24_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_71 = _mid_data_in_24_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_24_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_72 = _mid_data_in_24_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_24_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_73 = _mid_data_in_24_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_24_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_74 = _mid_data_in_24_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_24_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_75 = _mid_data_in_24_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_24_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_76 = _mid_data_in_24_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_24_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_77 = _mid_data_in_24_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_24_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_78 = _mid_data_in_24_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_24_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_79 = _mid_data_in_24_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_24_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_24_tdata_T_80 = _mid_data_in_24_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_24_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_66 = _mid_data_in_24_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_24_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_67 = _mid_data_in_24_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_24_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_68 = _mid_data_in_24_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_24_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_69 = _mid_data_in_24_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_24_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_70 = _mid_data_in_24_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_24_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_71 = _mid_data_in_24_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_24_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_72 = _mid_data_in_24_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_24_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_73 = _mid_data_in_24_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_24_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_74 = _mid_data_in_24_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_24_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_75 = _mid_data_in_24_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_24_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_76 = _mid_data_in_24_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_24_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_77 = _mid_data_in_24_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_24_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_78 = _mid_data_in_24_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_24_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_79 = _mid_data_in_24_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_24_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_24_tkeep_T_80 = _mid_data_in_24_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_24_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_97 = _T_100 < 32'h10 ? _mid_data_in_24_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_98 = _T_100 < 32'h10 & _mid_data_in_24_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_24_tdata = 32'h18 >= mid_count ? _GEN_97 : mid_m_axis_tdata[799:768]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_24_tkeep = 32'h18 >= mid_count ? _GEN_98 : mid_m_axis_tkeep[24]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_104 = 32'h19 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_25_tdata_T_3 = 32'h0 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_7 = 32'h1 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_11 = 32'h2 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_15 = 32'h3 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_19 = 32'h4 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_23 = 32'h5 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_27 = 32'h6 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_31 = 32'h7 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_35 = 32'h8 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_39 = 32'h9 == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_43 = 32'ha == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_47 = 32'hb == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_51 = 32'hc == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_55 = 32'hd == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_59 = 32'he == _T_104; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_25_tdata_T_63 = 32'hf == _T_104; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_25_tdata_T_65 = _mid_data_in_25_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_66 = _mid_data_in_25_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_25_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_67 = _mid_data_in_25_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_25_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_68 = _mid_data_in_25_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_25_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_69 = _mid_data_in_25_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_25_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_70 = _mid_data_in_25_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_25_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_71 = _mid_data_in_25_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_25_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_72 = _mid_data_in_25_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_25_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_73 = _mid_data_in_25_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_25_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_74 = _mid_data_in_25_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_25_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_75 = _mid_data_in_25_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_25_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_76 = _mid_data_in_25_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_25_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_77 = _mid_data_in_25_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_25_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_78 = _mid_data_in_25_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_25_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_79 = _mid_data_in_25_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_25_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_25_tdata_T_80 = _mid_data_in_25_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_25_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_66 = _mid_data_in_25_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_25_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_67 = _mid_data_in_25_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_25_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_68 = _mid_data_in_25_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_25_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_69 = _mid_data_in_25_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_25_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_70 = _mid_data_in_25_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_25_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_71 = _mid_data_in_25_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_25_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_72 = _mid_data_in_25_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_25_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_73 = _mid_data_in_25_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_25_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_74 = _mid_data_in_25_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_25_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_75 = _mid_data_in_25_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_25_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_76 = _mid_data_in_25_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_25_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_77 = _mid_data_in_25_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_25_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_78 = _mid_data_in_25_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_25_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_79 = _mid_data_in_25_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_25_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_25_tkeep_T_80 = _mid_data_in_25_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_25_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_101 = _T_104 < 32'h10 ? _mid_data_in_25_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_102 = _T_104 < 32'h10 & _mid_data_in_25_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_25_tdata = 32'h19 >= mid_count ? _GEN_101 : mid_m_axis_tdata[831:800]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_25_tkeep = 32'h19 >= mid_count ? _GEN_102 : mid_m_axis_tkeep[25]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_108 = 32'h1a - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_26_tdata_T_3 = 32'h0 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_7 = 32'h1 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_11 = 32'h2 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_15 = 32'h3 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_19 = 32'h4 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_23 = 32'h5 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_27 = 32'h6 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_31 = 32'h7 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_35 = 32'h8 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_39 = 32'h9 == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_43 = 32'ha == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_47 = 32'hb == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_51 = 32'hc == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_55 = 32'hd == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_59 = 32'he == _T_108; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_26_tdata_T_63 = 32'hf == _T_108; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_26_tdata_T_65 = _mid_data_in_26_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_66 = _mid_data_in_26_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_26_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_67 = _mid_data_in_26_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_26_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_68 = _mid_data_in_26_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_26_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_69 = _mid_data_in_26_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_26_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_70 = _mid_data_in_26_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_26_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_71 = _mid_data_in_26_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_26_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_72 = _mid_data_in_26_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_26_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_73 = _mid_data_in_26_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_26_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_74 = _mid_data_in_26_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_26_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_75 = _mid_data_in_26_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_26_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_76 = _mid_data_in_26_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_26_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_77 = _mid_data_in_26_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_26_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_78 = _mid_data_in_26_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_26_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_79 = _mid_data_in_26_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_26_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_26_tdata_T_80 = _mid_data_in_26_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_26_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_66 = _mid_data_in_26_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_26_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_67 = _mid_data_in_26_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_26_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_68 = _mid_data_in_26_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_26_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_69 = _mid_data_in_26_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_26_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_70 = _mid_data_in_26_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_26_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_71 = _mid_data_in_26_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_26_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_72 = _mid_data_in_26_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_26_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_73 = _mid_data_in_26_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_26_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_74 = _mid_data_in_26_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_26_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_75 = _mid_data_in_26_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_26_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_76 = _mid_data_in_26_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_26_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_77 = _mid_data_in_26_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_26_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_78 = _mid_data_in_26_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_26_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_79 = _mid_data_in_26_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_26_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_26_tkeep_T_80 = _mid_data_in_26_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_26_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_105 = _T_108 < 32'h10 ? _mid_data_in_26_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_106 = _T_108 < 32'h10 & _mid_data_in_26_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_26_tdata = 32'h1a >= mid_count ? _GEN_105 : mid_m_axis_tdata[863:832]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_26_tkeep = 32'h1a >= mid_count ? _GEN_106 : mid_m_axis_tkeep[26]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_112 = 32'h1b - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_27_tdata_T_3 = 32'h0 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_7 = 32'h1 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_11 = 32'h2 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_15 = 32'h3 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_19 = 32'h4 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_23 = 32'h5 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_27 = 32'h6 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_31 = 32'h7 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_35 = 32'h8 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_39 = 32'h9 == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_43 = 32'ha == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_47 = 32'hb == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_51 = 32'hc == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_55 = 32'hd == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_59 = 32'he == _T_112; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_27_tdata_T_63 = 32'hf == _T_112; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_27_tdata_T_65 = _mid_data_in_27_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_66 = _mid_data_in_27_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_27_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_67 = _mid_data_in_27_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_27_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_68 = _mid_data_in_27_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_27_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_69 = _mid_data_in_27_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_27_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_70 = _mid_data_in_27_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_27_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_71 = _mid_data_in_27_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_27_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_72 = _mid_data_in_27_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_27_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_73 = _mid_data_in_27_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_27_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_74 = _mid_data_in_27_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_27_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_75 = _mid_data_in_27_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_27_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_76 = _mid_data_in_27_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_27_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_77 = _mid_data_in_27_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_27_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_78 = _mid_data_in_27_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_27_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_79 = _mid_data_in_27_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_27_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_27_tdata_T_80 = _mid_data_in_27_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_27_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_66 = _mid_data_in_27_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_27_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_67 = _mid_data_in_27_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_27_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_68 = _mid_data_in_27_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_27_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_69 = _mid_data_in_27_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_27_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_70 = _mid_data_in_27_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_27_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_71 = _mid_data_in_27_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_27_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_72 = _mid_data_in_27_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_27_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_73 = _mid_data_in_27_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_27_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_74 = _mid_data_in_27_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_27_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_75 = _mid_data_in_27_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_27_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_76 = _mid_data_in_27_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_27_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_77 = _mid_data_in_27_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_27_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_78 = _mid_data_in_27_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_27_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_79 = _mid_data_in_27_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_27_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_27_tkeep_T_80 = _mid_data_in_27_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_27_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_109 = _T_112 < 32'h10 ? _mid_data_in_27_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_110 = _T_112 < 32'h10 & _mid_data_in_27_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_27_tdata = 32'h1b >= mid_count ? _GEN_109 : mid_m_axis_tdata[895:864]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_27_tkeep = 32'h1b >= mid_count ? _GEN_110 : mid_m_axis_tkeep[27]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_116 = 32'h1c - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_28_tdata_T_3 = 32'h0 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_7 = 32'h1 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_11 = 32'h2 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_15 = 32'h3 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_19 = 32'h4 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_23 = 32'h5 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_27 = 32'h6 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_31 = 32'h7 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_35 = 32'h8 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_39 = 32'h9 == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_43 = 32'ha == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_47 = 32'hb == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_51 = 32'hc == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_55 = 32'hd == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_59 = 32'he == _T_116; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_28_tdata_T_63 = 32'hf == _T_116; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_28_tdata_T_65 = _mid_data_in_28_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_66 = _mid_data_in_28_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_28_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_67 = _mid_data_in_28_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_28_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_68 = _mid_data_in_28_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_28_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_69 = _mid_data_in_28_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_28_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_70 = _mid_data_in_28_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_28_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_71 = _mid_data_in_28_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_28_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_72 = _mid_data_in_28_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_28_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_73 = _mid_data_in_28_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_28_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_74 = _mid_data_in_28_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_28_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_75 = _mid_data_in_28_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_28_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_76 = _mid_data_in_28_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_28_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_77 = _mid_data_in_28_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_28_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_78 = _mid_data_in_28_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_28_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_79 = _mid_data_in_28_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_28_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_28_tdata_T_80 = _mid_data_in_28_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_28_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_66 = _mid_data_in_28_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_28_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_67 = _mid_data_in_28_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_28_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_68 = _mid_data_in_28_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_28_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_69 = _mid_data_in_28_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_28_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_70 = _mid_data_in_28_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_28_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_71 = _mid_data_in_28_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_28_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_72 = _mid_data_in_28_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_28_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_73 = _mid_data_in_28_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_28_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_74 = _mid_data_in_28_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_28_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_75 = _mid_data_in_28_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_28_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_76 = _mid_data_in_28_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_28_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_77 = _mid_data_in_28_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_28_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_78 = _mid_data_in_28_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_28_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_79 = _mid_data_in_28_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_28_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_28_tkeep_T_80 = _mid_data_in_28_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_28_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_113 = _T_116 < 32'h10 ? _mid_data_in_28_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_114 = _T_116 < 32'h10 & _mid_data_in_28_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_28_tdata = 32'h1c >= mid_count ? _GEN_113 : mid_m_axis_tdata[927:896]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_28_tkeep = 32'h1c >= mid_count ? _GEN_114 : mid_m_axis_tkeep[28]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_120 = 32'h1d - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_29_tdata_T_3 = 32'h0 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_7 = 32'h1 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_11 = 32'h2 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_15 = 32'h3 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_19 = 32'h4 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_23 = 32'h5 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_27 = 32'h6 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_31 = 32'h7 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_35 = 32'h8 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_39 = 32'h9 == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_43 = 32'ha == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_47 = 32'hb == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_51 = 32'hc == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_55 = 32'hd == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_59 = 32'he == _T_120; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_29_tdata_T_63 = 32'hf == _T_120; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_29_tdata_T_65 = _mid_data_in_29_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_66 = _mid_data_in_29_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_29_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_67 = _mid_data_in_29_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_29_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_68 = _mid_data_in_29_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_29_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_69 = _mid_data_in_29_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_29_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_70 = _mid_data_in_29_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_29_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_71 = _mid_data_in_29_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_29_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_72 = _mid_data_in_29_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_29_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_73 = _mid_data_in_29_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_29_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_74 = _mid_data_in_29_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_29_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_75 = _mid_data_in_29_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_29_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_76 = _mid_data_in_29_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_29_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_77 = _mid_data_in_29_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_29_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_78 = _mid_data_in_29_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_29_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_79 = _mid_data_in_29_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_29_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_29_tdata_T_80 = _mid_data_in_29_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_29_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_66 = _mid_data_in_29_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_29_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_67 = _mid_data_in_29_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_29_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_68 = _mid_data_in_29_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_29_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_69 = _mid_data_in_29_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_29_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_70 = _mid_data_in_29_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_29_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_71 = _mid_data_in_29_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_29_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_72 = _mid_data_in_29_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_29_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_73 = _mid_data_in_29_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_29_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_74 = _mid_data_in_29_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_29_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_75 = _mid_data_in_29_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_29_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_76 = _mid_data_in_29_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_29_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_77 = _mid_data_in_29_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_29_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_78 = _mid_data_in_29_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_29_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_79 = _mid_data_in_29_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_29_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_29_tkeep_T_80 = _mid_data_in_29_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_29_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_117 = _T_120 < 32'h10 ? _mid_data_in_29_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_118 = _T_120 < 32'h10 & _mid_data_in_29_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_29_tdata = 32'h1d >= mid_count ? _GEN_117 : mid_m_axis_tdata[959:928]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_29_tkeep = 32'h1d >= mid_count ? _GEN_118 : mid_m_axis_tkeep[29]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_124 = 32'h1e - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_30_tdata_T_3 = 32'h0 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_7 = 32'h1 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_11 = 32'h2 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_15 = 32'h3 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_19 = 32'h4 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_23 = 32'h5 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_27 = 32'h6 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_31 = 32'h7 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_35 = 32'h8 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_39 = 32'h9 == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_43 = 32'ha == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_47 = 32'hb == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_51 = 32'hc == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_55 = 32'hd == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_59 = 32'he == _T_124; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_30_tdata_T_63 = 32'hf == _T_124; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_30_tdata_T_65 = _mid_data_in_30_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_66 = _mid_data_in_30_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_30_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_67 = _mid_data_in_30_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_30_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_68 = _mid_data_in_30_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_30_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_69 = _mid_data_in_30_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_30_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_70 = _mid_data_in_30_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_30_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_71 = _mid_data_in_30_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_30_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_72 = _mid_data_in_30_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_30_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_73 = _mid_data_in_30_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_30_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_74 = _mid_data_in_30_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_30_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_75 = _mid_data_in_30_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_30_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_76 = _mid_data_in_30_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_30_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_77 = _mid_data_in_30_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_30_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_78 = _mid_data_in_30_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_30_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_79 = _mid_data_in_30_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_30_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_30_tdata_T_80 = _mid_data_in_30_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_30_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_66 = _mid_data_in_30_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_30_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_67 = _mid_data_in_30_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_30_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_68 = _mid_data_in_30_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_30_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_69 = _mid_data_in_30_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_30_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_70 = _mid_data_in_30_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_30_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_71 = _mid_data_in_30_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_30_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_72 = _mid_data_in_30_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_30_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_73 = _mid_data_in_30_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_30_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_74 = _mid_data_in_30_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_30_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_75 = _mid_data_in_30_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_30_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_76 = _mid_data_in_30_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_30_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_77 = _mid_data_in_30_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_30_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_78 = _mid_data_in_30_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_30_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_79 = _mid_data_in_30_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_30_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_30_tkeep_T_80 = _mid_data_in_30_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_30_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_121 = _T_124 < 32'h10 ? _mid_data_in_30_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_122 = _T_124 < 32'h10 & _mid_data_in_30_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_30_tdata = 32'h1e >= mid_count ? _GEN_121 : mid_m_axis_tdata[991:960]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_30_tkeep = 32'h1e >= mid_count ? _GEN_122 : mid_m_axis_tkeep[30]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_128 = 32'h1f - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_31_tdata_T_3 = 32'h0 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_7 = 32'h1 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_11 = 32'h2 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_15 = 32'h3 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_19 = 32'h4 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_23 = 32'h5 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_27 = 32'h6 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_31 = 32'h7 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_35 = 32'h8 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_39 = 32'h9 == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_43 = 32'ha == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_47 = 32'hb == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_51 = 32'hc == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_55 = 32'hd == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_59 = 32'he == _T_128; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_31_tdata_T_63 = 32'hf == _T_128; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_31_tdata_T_65 = _mid_data_in_31_tdata_T_63 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_66 = _mid_data_in_31_tdata_T_59 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_31_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_67 = _mid_data_in_31_tdata_T_55 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_31_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_68 = _mid_data_in_31_tdata_T_51 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_31_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_69 = _mid_data_in_31_tdata_T_47 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_31_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_70 = _mid_data_in_31_tdata_T_43 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_31_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_71 = _mid_data_in_31_tdata_T_39 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_31_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_72 = _mid_data_in_31_tdata_T_35 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_31_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_73 = _mid_data_in_31_tdata_T_31 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_31_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_74 = _mid_data_in_31_tdata_T_27 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_31_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_75 = _mid_data_in_31_tdata_T_23 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_31_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_76 = _mid_data_in_31_tdata_T_19 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_31_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_77 = _mid_data_in_31_tdata_T_15 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_31_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_78 = _mid_data_in_31_tdata_T_11 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_31_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_79 = _mid_data_in_31_tdata_T_7 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_31_tdata_T_78; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_31_tdata_T_80 = _mid_data_in_31_tdata_T_3 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_31_tdata_T_79; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_66 = _mid_data_in_31_tdata_T_59 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_31_tdata_T_63 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_67 = _mid_data_in_31_tdata_T_55 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_31_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_68 = _mid_data_in_31_tdata_T_51 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_31_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_69 = _mid_data_in_31_tdata_T_47 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_31_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_70 = _mid_data_in_31_tdata_T_43 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_31_tkeep_T_69; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_71 = _mid_data_in_31_tdata_T_39 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_31_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_72 = _mid_data_in_31_tdata_T_35 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_31_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_73 = _mid_data_in_31_tdata_T_31 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_31_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_74 = _mid_data_in_31_tdata_T_27 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_31_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_75 = _mid_data_in_31_tdata_T_23 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_31_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_76 = _mid_data_in_31_tdata_T_19 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_31_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_77 = _mid_data_in_31_tdata_T_15 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_31_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_78 = _mid_data_in_31_tdata_T_11 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_31_tkeep_T_77
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_79 = _mid_data_in_31_tdata_T_7 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_31_tkeep_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_31_tkeep_T_80 = _mid_data_in_31_tdata_T_3 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_31_tkeep_T_79; // @[Mux.scala 98:16]
  wire [31:0] _GEN_125 = _T_128 < 32'h10 ? _mid_data_in_31_tdata_T_80 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_126 = _T_128 < 32'h10 & _mid_data_in_31_tkeep_T_80; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_31_tdata = 32'h1f >= mid_count ? _GEN_125 : mid_m_axis_tdata[1023:992]; // @[bfs_remote.scala 70:29 bfs_remote.scala 64:17]
  wire  mid_data_in_31_tkeep = 32'h1f >= mid_count ? _GEN_126 : mid_m_axis_tkeep[31]; // @[bfs_remote.scala 70:29 bfs_remote.scala 65:17]
  wire [31:0] _T_132 = 32'h20 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_32_tdata_T_2 = 32'h0 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_6 = 32'h1 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_10 = 32'h2 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_14 = 32'h3 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_18 = 32'h4 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_22 = 32'h5 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_26 = 32'h6 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_30 = 32'h7 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_34 = 32'h8 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_38 = 32'h9 == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_42 = 32'ha == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_46 = 32'hb == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_50 = 32'hc == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_54 = 32'hd == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_58 = 32'he == _T_132; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_32_tdata_T_62 = 32'hf == _T_132; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_32_tdata_T_64 = _mid_data_in_32_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_65 = _mid_data_in_32_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_32_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_66 = _mid_data_in_32_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_32_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_67 = _mid_data_in_32_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_32_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_68 = _mid_data_in_32_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_32_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_69 = _mid_data_in_32_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_32_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_70 = _mid_data_in_32_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_32_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_71 = _mid_data_in_32_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_32_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_72 = _mid_data_in_32_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_32_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_73 = _mid_data_in_32_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_32_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_74 = _mid_data_in_32_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_32_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_75 = _mid_data_in_32_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_32_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_76 = _mid_data_in_32_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_32_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_77 = _mid_data_in_32_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_32_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_78 = _mid_data_in_32_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_32_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_32_tdata_T_79 = _mid_data_in_32_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_32_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_65 = _mid_data_in_32_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_32_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_66 = _mid_data_in_32_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_32_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_67 = _mid_data_in_32_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_32_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_68 = _mid_data_in_32_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_32_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_69 = _mid_data_in_32_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_32_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_70 = _mid_data_in_32_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_32_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_71 = _mid_data_in_32_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_32_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_72 = _mid_data_in_32_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_32_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_73 = _mid_data_in_32_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_32_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_74 = _mid_data_in_32_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_32_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_75 = _mid_data_in_32_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_32_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_76 = _mid_data_in_32_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_32_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_77 = _mid_data_in_32_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_32_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_78 = _mid_data_in_32_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_32_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_32_tkeep_T_79 = _mid_data_in_32_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_32_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_129 = _T_132 < 32'h10 ? _mid_data_in_32_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_130 = _T_132 < 32'h10 & _mid_data_in_32_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_32_tdata = 32'h20 >= mid_count ? _GEN_129 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_32_tkeep = 32'h20 >= mid_count & _GEN_130; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_136 = 32'h21 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_33_tdata_T_2 = 32'h0 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_6 = 32'h1 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_10 = 32'h2 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_14 = 32'h3 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_18 = 32'h4 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_22 = 32'h5 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_26 = 32'h6 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_30 = 32'h7 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_34 = 32'h8 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_38 = 32'h9 == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_42 = 32'ha == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_46 = 32'hb == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_50 = 32'hc == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_54 = 32'hd == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_58 = 32'he == _T_136; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_33_tdata_T_62 = 32'hf == _T_136; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_33_tdata_T_64 = _mid_data_in_33_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_65 = _mid_data_in_33_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_33_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_66 = _mid_data_in_33_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_33_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_67 = _mid_data_in_33_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_33_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_68 = _mid_data_in_33_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_33_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_69 = _mid_data_in_33_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_33_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_70 = _mid_data_in_33_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_33_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_71 = _mid_data_in_33_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_33_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_72 = _mid_data_in_33_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_33_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_73 = _mid_data_in_33_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_33_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_74 = _mid_data_in_33_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_33_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_75 = _mid_data_in_33_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_33_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_76 = _mid_data_in_33_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_33_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_77 = _mid_data_in_33_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_33_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_78 = _mid_data_in_33_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_33_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_33_tdata_T_79 = _mid_data_in_33_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_33_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_65 = _mid_data_in_33_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_33_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_66 = _mid_data_in_33_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_33_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_67 = _mid_data_in_33_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_33_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_68 = _mid_data_in_33_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_33_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_69 = _mid_data_in_33_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_33_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_70 = _mid_data_in_33_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_33_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_71 = _mid_data_in_33_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_33_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_72 = _mid_data_in_33_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_33_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_73 = _mid_data_in_33_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_33_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_74 = _mid_data_in_33_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_33_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_75 = _mid_data_in_33_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_33_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_76 = _mid_data_in_33_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_33_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_77 = _mid_data_in_33_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_33_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_78 = _mid_data_in_33_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_33_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_33_tkeep_T_79 = _mid_data_in_33_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_33_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_133 = _T_136 < 32'h10 ? _mid_data_in_33_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_134 = _T_136 < 32'h10 & _mid_data_in_33_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_33_tdata = 32'h21 >= mid_count ? _GEN_133 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_33_tkeep = 32'h21 >= mid_count & _GEN_134; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_140 = 32'h22 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_34_tdata_T_2 = 32'h0 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_6 = 32'h1 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_10 = 32'h2 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_14 = 32'h3 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_18 = 32'h4 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_22 = 32'h5 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_26 = 32'h6 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_30 = 32'h7 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_34 = 32'h8 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_38 = 32'h9 == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_42 = 32'ha == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_46 = 32'hb == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_50 = 32'hc == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_54 = 32'hd == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_58 = 32'he == _T_140; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_34_tdata_T_62 = 32'hf == _T_140; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_34_tdata_T_64 = _mid_data_in_34_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_65 = _mid_data_in_34_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_34_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_66 = _mid_data_in_34_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_34_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_67 = _mid_data_in_34_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_34_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_68 = _mid_data_in_34_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_34_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_69 = _mid_data_in_34_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_34_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_70 = _mid_data_in_34_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_34_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_71 = _mid_data_in_34_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_34_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_72 = _mid_data_in_34_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_34_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_73 = _mid_data_in_34_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_34_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_74 = _mid_data_in_34_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_34_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_75 = _mid_data_in_34_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_34_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_76 = _mid_data_in_34_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_34_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_77 = _mid_data_in_34_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_34_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_78 = _mid_data_in_34_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_34_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_34_tdata_T_79 = _mid_data_in_34_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_34_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_65 = _mid_data_in_34_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_34_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_66 = _mid_data_in_34_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_34_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_67 = _mid_data_in_34_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_34_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_68 = _mid_data_in_34_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_34_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_69 = _mid_data_in_34_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_34_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_70 = _mid_data_in_34_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_34_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_71 = _mid_data_in_34_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_34_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_72 = _mid_data_in_34_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_34_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_73 = _mid_data_in_34_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_34_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_74 = _mid_data_in_34_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_34_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_75 = _mid_data_in_34_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_34_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_76 = _mid_data_in_34_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_34_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_77 = _mid_data_in_34_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_34_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_78 = _mid_data_in_34_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_34_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_34_tkeep_T_79 = _mid_data_in_34_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_34_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_137 = _T_140 < 32'h10 ? _mid_data_in_34_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_138 = _T_140 < 32'h10 & _mid_data_in_34_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_34_tdata = 32'h22 >= mid_count ? _GEN_137 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_34_tkeep = 32'h22 >= mid_count & _GEN_138; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_144 = 32'h23 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_35_tdata_T_2 = 32'h0 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_6 = 32'h1 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_10 = 32'h2 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_14 = 32'h3 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_18 = 32'h4 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_22 = 32'h5 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_26 = 32'h6 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_30 = 32'h7 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_34 = 32'h8 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_38 = 32'h9 == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_42 = 32'ha == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_46 = 32'hb == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_50 = 32'hc == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_54 = 32'hd == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_58 = 32'he == _T_144; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_35_tdata_T_62 = 32'hf == _T_144; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_35_tdata_T_64 = _mid_data_in_35_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_65 = _mid_data_in_35_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_35_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_66 = _mid_data_in_35_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_35_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_67 = _mid_data_in_35_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_35_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_68 = _mid_data_in_35_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_35_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_69 = _mid_data_in_35_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_35_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_70 = _mid_data_in_35_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_35_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_71 = _mid_data_in_35_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_35_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_72 = _mid_data_in_35_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_35_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_73 = _mid_data_in_35_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_35_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_74 = _mid_data_in_35_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_35_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_75 = _mid_data_in_35_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_35_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_76 = _mid_data_in_35_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_35_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_77 = _mid_data_in_35_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_35_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_78 = _mid_data_in_35_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_35_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_35_tdata_T_79 = _mid_data_in_35_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_35_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_65 = _mid_data_in_35_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_35_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_66 = _mid_data_in_35_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_35_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_67 = _mid_data_in_35_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_35_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_68 = _mid_data_in_35_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_35_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_69 = _mid_data_in_35_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_35_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_70 = _mid_data_in_35_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_35_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_71 = _mid_data_in_35_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_35_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_72 = _mid_data_in_35_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_35_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_73 = _mid_data_in_35_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_35_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_74 = _mid_data_in_35_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_35_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_75 = _mid_data_in_35_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_35_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_76 = _mid_data_in_35_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_35_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_77 = _mid_data_in_35_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_35_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_78 = _mid_data_in_35_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_35_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_35_tkeep_T_79 = _mid_data_in_35_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_35_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_141 = _T_144 < 32'h10 ? _mid_data_in_35_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_142 = _T_144 < 32'h10 & _mid_data_in_35_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_35_tdata = 32'h23 >= mid_count ? _GEN_141 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_35_tkeep = 32'h23 >= mid_count & _GEN_142; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_148 = 32'h24 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_36_tdata_T_2 = 32'h0 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_6 = 32'h1 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_10 = 32'h2 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_14 = 32'h3 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_18 = 32'h4 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_22 = 32'h5 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_26 = 32'h6 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_30 = 32'h7 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_34 = 32'h8 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_38 = 32'h9 == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_42 = 32'ha == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_46 = 32'hb == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_50 = 32'hc == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_54 = 32'hd == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_58 = 32'he == _T_148; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_36_tdata_T_62 = 32'hf == _T_148; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_36_tdata_T_64 = _mid_data_in_36_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_65 = _mid_data_in_36_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_36_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_66 = _mid_data_in_36_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_36_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_67 = _mid_data_in_36_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_36_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_68 = _mid_data_in_36_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_36_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_69 = _mid_data_in_36_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_36_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_70 = _mid_data_in_36_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_36_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_71 = _mid_data_in_36_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_36_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_72 = _mid_data_in_36_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_36_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_73 = _mid_data_in_36_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_36_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_74 = _mid_data_in_36_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_36_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_75 = _mid_data_in_36_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_36_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_76 = _mid_data_in_36_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_36_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_77 = _mid_data_in_36_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_36_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_78 = _mid_data_in_36_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_36_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_36_tdata_T_79 = _mid_data_in_36_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_36_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_65 = _mid_data_in_36_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_36_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_66 = _mid_data_in_36_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_36_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_67 = _mid_data_in_36_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_36_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_68 = _mid_data_in_36_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_36_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_69 = _mid_data_in_36_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_36_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_70 = _mid_data_in_36_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_36_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_71 = _mid_data_in_36_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_36_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_72 = _mid_data_in_36_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_36_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_73 = _mid_data_in_36_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_36_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_74 = _mid_data_in_36_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_36_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_75 = _mid_data_in_36_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_36_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_76 = _mid_data_in_36_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_36_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_77 = _mid_data_in_36_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_36_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_78 = _mid_data_in_36_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_36_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_36_tkeep_T_79 = _mid_data_in_36_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_36_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_145 = _T_148 < 32'h10 ? _mid_data_in_36_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_146 = _T_148 < 32'h10 & _mid_data_in_36_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_36_tdata = 32'h24 >= mid_count ? _GEN_145 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_36_tkeep = 32'h24 >= mid_count & _GEN_146; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_152 = 32'h25 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_37_tdata_T_2 = 32'h0 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_6 = 32'h1 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_10 = 32'h2 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_14 = 32'h3 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_18 = 32'h4 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_22 = 32'h5 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_26 = 32'h6 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_30 = 32'h7 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_34 = 32'h8 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_38 = 32'h9 == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_42 = 32'ha == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_46 = 32'hb == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_50 = 32'hc == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_54 = 32'hd == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_58 = 32'he == _T_152; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_37_tdata_T_62 = 32'hf == _T_152; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_37_tdata_T_64 = _mid_data_in_37_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_65 = _mid_data_in_37_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_37_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_66 = _mid_data_in_37_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_37_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_67 = _mid_data_in_37_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_37_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_68 = _mid_data_in_37_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_37_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_69 = _mid_data_in_37_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_37_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_70 = _mid_data_in_37_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_37_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_71 = _mid_data_in_37_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_37_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_72 = _mid_data_in_37_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_37_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_73 = _mid_data_in_37_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_37_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_74 = _mid_data_in_37_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_37_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_75 = _mid_data_in_37_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_37_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_76 = _mid_data_in_37_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_37_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_77 = _mid_data_in_37_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_37_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_78 = _mid_data_in_37_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_37_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_37_tdata_T_79 = _mid_data_in_37_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_37_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_65 = _mid_data_in_37_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_37_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_66 = _mid_data_in_37_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_37_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_67 = _mid_data_in_37_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_37_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_68 = _mid_data_in_37_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_37_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_69 = _mid_data_in_37_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_37_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_70 = _mid_data_in_37_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_37_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_71 = _mid_data_in_37_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_37_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_72 = _mid_data_in_37_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_37_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_73 = _mid_data_in_37_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_37_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_74 = _mid_data_in_37_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_37_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_75 = _mid_data_in_37_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_37_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_76 = _mid_data_in_37_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_37_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_77 = _mid_data_in_37_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_37_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_78 = _mid_data_in_37_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_37_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_37_tkeep_T_79 = _mid_data_in_37_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_37_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_149 = _T_152 < 32'h10 ? _mid_data_in_37_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_150 = _T_152 < 32'h10 & _mid_data_in_37_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_37_tdata = 32'h25 >= mid_count ? _GEN_149 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_37_tkeep = 32'h25 >= mid_count & _GEN_150; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_156 = 32'h26 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_38_tdata_T_2 = 32'h0 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_6 = 32'h1 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_10 = 32'h2 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_14 = 32'h3 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_18 = 32'h4 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_22 = 32'h5 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_26 = 32'h6 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_30 = 32'h7 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_34 = 32'h8 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_38 = 32'h9 == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_42 = 32'ha == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_46 = 32'hb == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_50 = 32'hc == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_54 = 32'hd == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_58 = 32'he == _T_156; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_38_tdata_T_62 = 32'hf == _T_156; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_38_tdata_T_64 = _mid_data_in_38_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_65 = _mid_data_in_38_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_38_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_66 = _mid_data_in_38_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_38_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_67 = _mid_data_in_38_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_38_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_68 = _mid_data_in_38_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_38_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_69 = _mid_data_in_38_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_38_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_70 = _mid_data_in_38_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_38_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_71 = _mid_data_in_38_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_38_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_72 = _mid_data_in_38_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_38_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_73 = _mid_data_in_38_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_38_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_74 = _mid_data_in_38_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_38_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_75 = _mid_data_in_38_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_38_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_76 = _mid_data_in_38_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_38_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_77 = _mid_data_in_38_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_38_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_78 = _mid_data_in_38_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_38_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_38_tdata_T_79 = _mid_data_in_38_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_38_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_65 = _mid_data_in_38_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_38_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_66 = _mid_data_in_38_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_38_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_67 = _mid_data_in_38_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_38_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_68 = _mid_data_in_38_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_38_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_69 = _mid_data_in_38_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_38_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_70 = _mid_data_in_38_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_38_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_71 = _mid_data_in_38_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_38_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_72 = _mid_data_in_38_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_38_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_73 = _mid_data_in_38_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_38_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_74 = _mid_data_in_38_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_38_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_75 = _mid_data_in_38_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_38_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_76 = _mid_data_in_38_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_38_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_77 = _mid_data_in_38_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_38_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_78 = _mid_data_in_38_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_38_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_38_tkeep_T_79 = _mid_data_in_38_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_38_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_153 = _T_156 < 32'h10 ? _mid_data_in_38_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_154 = _T_156 < 32'h10 & _mid_data_in_38_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_38_tdata = 32'h26 >= mid_count ? _GEN_153 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_38_tkeep = 32'h26 >= mid_count & _GEN_154; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_160 = 32'h27 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_39_tdata_T_2 = 32'h0 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_6 = 32'h1 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_10 = 32'h2 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_14 = 32'h3 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_18 = 32'h4 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_22 = 32'h5 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_26 = 32'h6 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_30 = 32'h7 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_34 = 32'h8 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_38 = 32'h9 == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_42 = 32'ha == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_46 = 32'hb == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_50 = 32'hc == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_54 = 32'hd == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_58 = 32'he == _T_160; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_39_tdata_T_62 = 32'hf == _T_160; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_39_tdata_T_64 = _mid_data_in_39_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_65 = _mid_data_in_39_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_39_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_66 = _mid_data_in_39_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_39_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_67 = _mid_data_in_39_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_39_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_68 = _mid_data_in_39_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_39_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_69 = _mid_data_in_39_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_39_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_70 = _mid_data_in_39_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_39_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_71 = _mid_data_in_39_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_39_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_72 = _mid_data_in_39_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_39_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_73 = _mid_data_in_39_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_39_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_74 = _mid_data_in_39_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_39_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_75 = _mid_data_in_39_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_39_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_76 = _mid_data_in_39_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_39_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_77 = _mid_data_in_39_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_39_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_78 = _mid_data_in_39_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_39_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_39_tdata_T_79 = _mid_data_in_39_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_39_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_65 = _mid_data_in_39_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_39_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_66 = _mid_data_in_39_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_39_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_67 = _mid_data_in_39_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_39_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_68 = _mid_data_in_39_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_39_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_69 = _mid_data_in_39_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_39_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_70 = _mid_data_in_39_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_39_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_71 = _mid_data_in_39_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_39_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_72 = _mid_data_in_39_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_39_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_73 = _mid_data_in_39_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_39_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_74 = _mid_data_in_39_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_39_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_75 = _mid_data_in_39_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_39_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_76 = _mid_data_in_39_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_39_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_77 = _mid_data_in_39_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_39_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_78 = _mid_data_in_39_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_39_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_39_tkeep_T_79 = _mid_data_in_39_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_39_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_157 = _T_160 < 32'h10 ? _mid_data_in_39_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_158 = _T_160 < 32'h10 & _mid_data_in_39_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_39_tdata = 32'h27 >= mid_count ? _GEN_157 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_39_tkeep = 32'h27 >= mid_count & _GEN_158; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_164 = 32'h28 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_40_tdata_T_2 = 32'h0 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_6 = 32'h1 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_10 = 32'h2 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_14 = 32'h3 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_18 = 32'h4 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_22 = 32'h5 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_26 = 32'h6 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_30 = 32'h7 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_34 = 32'h8 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_38 = 32'h9 == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_42 = 32'ha == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_46 = 32'hb == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_50 = 32'hc == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_54 = 32'hd == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_58 = 32'he == _T_164; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_40_tdata_T_62 = 32'hf == _T_164; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_40_tdata_T_64 = _mid_data_in_40_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_65 = _mid_data_in_40_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_40_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_66 = _mid_data_in_40_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_40_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_67 = _mid_data_in_40_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_40_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_68 = _mid_data_in_40_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_40_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_69 = _mid_data_in_40_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_40_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_70 = _mid_data_in_40_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_40_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_71 = _mid_data_in_40_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_40_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_72 = _mid_data_in_40_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_40_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_73 = _mid_data_in_40_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_40_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_74 = _mid_data_in_40_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_40_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_75 = _mid_data_in_40_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_40_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_76 = _mid_data_in_40_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_40_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_77 = _mid_data_in_40_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_40_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_78 = _mid_data_in_40_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_40_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_40_tdata_T_79 = _mid_data_in_40_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_40_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_65 = _mid_data_in_40_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_40_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_66 = _mid_data_in_40_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_40_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_67 = _mid_data_in_40_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_40_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_68 = _mid_data_in_40_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_40_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_69 = _mid_data_in_40_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_40_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_70 = _mid_data_in_40_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_40_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_71 = _mid_data_in_40_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_40_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_72 = _mid_data_in_40_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_40_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_73 = _mid_data_in_40_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_40_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_74 = _mid_data_in_40_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_40_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_75 = _mid_data_in_40_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_40_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_76 = _mid_data_in_40_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_40_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_77 = _mid_data_in_40_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_40_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_78 = _mid_data_in_40_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_40_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_40_tkeep_T_79 = _mid_data_in_40_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_40_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_161 = _T_164 < 32'h10 ? _mid_data_in_40_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_162 = _T_164 < 32'h10 & _mid_data_in_40_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_40_tdata = 32'h28 >= mid_count ? _GEN_161 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_40_tkeep = 32'h28 >= mid_count & _GEN_162; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_168 = 32'h29 - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_41_tdata_T_2 = 32'h0 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_6 = 32'h1 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_10 = 32'h2 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_14 = 32'h3 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_18 = 32'h4 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_22 = 32'h5 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_26 = 32'h6 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_30 = 32'h7 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_34 = 32'h8 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_38 = 32'h9 == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_42 = 32'ha == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_46 = 32'hb == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_50 = 32'hc == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_54 = 32'hd == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_58 = 32'he == _T_168; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_41_tdata_T_62 = 32'hf == _T_168; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_41_tdata_T_64 = _mid_data_in_41_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_65 = _mid_data_in_41_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_41_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_66 = _mid_data_in_41_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_41_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_67 = _mid_data_in_41_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_41_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_68 = _mid_data_in_41_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_41_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_69 = _mid_data_in_41_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_41_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_70 = _mid_data_in_41_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_41_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_71 = _mid_data_in_41_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_41_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_72 = _mid_data_in_41_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_41_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_73 = _mid_data_in_41_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_41_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_74 = _mid_data_in_41_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_41_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_75 = _mid_data_in_41_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_41_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_76 = _mid_data_in_41_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_41_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_77 = _mid_data_in_41_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_41_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_78 = _mid_data_in_41_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_41_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_41_tdata_T_79 = _mid_data_in_41_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_41_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_65 = _mid_data_in_41_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_41_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_66 = _mid_data_in_41_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_41_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_67 = _mid_data_in_41_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_41_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_68 = _mid_data_in_41_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_41_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_69 = _mid_data_in_41_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_41_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_70 = _mid_data_in_41_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_41_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_71 = _mid_data_in_41_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_41_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_72 = _mid_data_in_41_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_41_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_73 = _mid_data_in_41_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_41_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_74 = _mid_data_in_41_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_41_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_75 = _mid_data_in_41_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_41_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_76 = _mid_data_in_41_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_41_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_77 = _mid_data_in_41_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_41_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_78 = _mid_data_in_41_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_41_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_41_tkeep_T_79 = _mid_data_in_41_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_41_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_165 = _T_168 < 32'h10 ? _mid_data_in_41_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_166 = _T_168 < 32'h10 & _mid_data_in_41_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_41_tdata = 32'h29 >= mid_count ? _GEN_165 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_41_tkeep = 32'h29 >= mid_count & _GEN_166; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_172 = 32'h2a - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_42_tdata_T_2 = 32'h0 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_6 = 32'h1 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_10 = 32'h2 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_14 = 32'h3 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_18 = 32'h4 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_22 = 32'h5 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_26 = 32'h6 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_30 = 32'h7 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_34 = 32'h8 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_38 = 32'h9 == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_42 = 32'ha == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_46 = 32'hb == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_50 = 32'hc == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_54 = 32'hd == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_58 = 32'he == _T_172; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_42_tdata_T_62 = 32'hf == _T_172; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_42_tdata_T_64 = _mid_data_in_42_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_65 = _mid_data_in_42_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_42_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_66 = _mid_data_in_42_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_42_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_67 = _mid_data_in_42_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_42_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_68 = _mid_data_in_42_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_42_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_69 = _mid_data_in_42_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_42_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_70 = _mid_data_in_42_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_42_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_71 = _mid_data_in_42_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_42_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_72 = _mid_data_in_42_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_42_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_73 = _mid_data_in_42_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_42_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_74 = _mid_data_in_42_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_42_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_75 = _mid_data_in_42_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_42_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_76 = _mid_data_in_42_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_42_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_77 = _mid_data_in_42_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_42_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_78 = _mid_data_in_42_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_42_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_42_tdata_T_79 = _mid_data_in_42_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_42_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_65 = _mid_data_in_42_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_42_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_66 = _mid_data_in_42_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_42_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_67 = _mid_data_in_42_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_42_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_68 = _mid_data_in_42_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_42_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_69 = _mid_data_in_42_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_42_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_70 = _mid_data_in_42_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_42_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_71 = _mid_data_in_42_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_42_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_72 = _mid_data_in_42_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_42_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_73 = _mid_data_in_42_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_42_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_74 = _mid_data_in_42_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_42_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_75 = _mid_data_in_42_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_42_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_76 = _mid_data_in_42_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_42_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_77 = _mid_data_in_42_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_42_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_78 = _mid_data_in_42_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_42_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_42_tkeep_T_79 = _mid_data_in_42_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_42_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_169 = _T_172 < 32'h10 ? _mid_data_in_42_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_170 = _T_172 < 32'h10 & _mid_data_in_42_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_42_tdata = 32'h2a >= mid_count ? _GEN_169 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_42_tkeep = 32'h2a >= mid_count & _GEN_170; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_176 = 32'h2b - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_43_tdata_T_2 = 32'h0 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_6 = 32'h1 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_10 = 32'h2 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_14 = 32'h3 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_18 = 32'h4 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_22 = 32'h5 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_26 = 32'h6 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_30 = 32'h7 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_34 = 32'h8 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_38 = 32'h9 == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_42 = 32'ha == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_46 = 32'hb == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_50 = 32'hc == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_54 = 32'hd == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_58 = 32'he == _T_176; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_43_tdata_T_62 = 32'hf == _T_176; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_43_tdata_T_64 = _mid_data_in_43_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_65 = _mid_data_in_43_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_43_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_66 = _mid_data_in_43_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_43_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_67 = _mid_data_in_43_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_43_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_68 = _mid_data_in_43_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_43_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_69 = _mid_data_in_43_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_43_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_70 = _mid_data_in_43_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_43_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_71 = _mid_data_in_43_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_43_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_72 = _mid_data_in_43_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_43_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_73 = _mid_data_in_43_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_43_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_74 = _mid_data_in_43_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_43_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_75 = _mid_data_in_43_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_43_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_76 = _mid_data_in_43_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_43_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_77 = _mid_data_in_43_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_43_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_78 = _mid_data_in_43_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_43_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_43_tdata_T_79 = _mid_data_in_43_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_43_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_65 = _mid_data_in_43_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_43_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_66 = _mid_data_in_43_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_43_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_67 = _mid_data_in_43_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_43_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_68 = _mid_data_in_43_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_43_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_69 = _mid_data_in_43_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_43_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_70 = _mid_data_in_43_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_43_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_71 = _mid_data_in_43_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_43_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_72 = _mid_data_in_43_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_43_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_73 = _mid_data_in_43_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_43_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_74 = _mid_data_in_43_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_43_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_75 = _mid_data_in_43_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_43_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_76 = _mid_data_in_43_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_43_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_77 = _mid_data_in_43_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_43_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_78 = _mid_data_in_43_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_43_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_43_tkeep_T_79 = _mid_data_in_43_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_43_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_173 = _T_176 < 32'h10 ? _mid_data_in_43_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_174 = _T_176 < 32'h10 & _mid_data_in_43_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_43_tdata = 32'h2b >= mid_count ? _GEN_173 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_43_tkeep = 32'h2b >= mid_count & _GEN_174; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_180 = 32'h2c - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_44_tdata_T_2 = 32'h0 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_6 = 32'h1 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_10 = 32'h2 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_14 = 32'h3 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_18 = 32'h4 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_22 = 32'h5 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_26 = 32'h6 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_30 = 32'h7 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_34 = 32'h8 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_38 = 32'h9 == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_42 = 32'ha == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_46 = 32'hb == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_50 = 32'hc == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_54 = 32'hd == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_58 = 32'he == _T_180; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_44_tdata_T_62 = 32'hf == _T_180; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_44_tdata_T_64 = _mid_data_in_44_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_65 = _mid_data_in_44_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_44_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_66 = _mid_data_in_44_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_44_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_67 = _mid_data_in_44_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_44_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_68 = _mid_data_in_44_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_44_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_69 = _mid_data_in_44_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_44_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_70 = _mid_data_in_44_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_44_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_71 = _mid_data_in_44_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_44_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_72 = _mid_data_in_44_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_44_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_73 = _mid_data_in_44_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_44_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_74 = _mid_data_in_44_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_44_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_75 = _mid_data_in_44_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_44_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_76 = _mid_data_in_44_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_44_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_77 = _mid_data_in_44_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_44_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_78 = _mid_data_in_44_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_44_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_44_tdata_T_79 = _mid_data_in_44_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_44_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_65 = _mid_data_in_44_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_44_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_66 = _mid_data_in_44_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_44_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_67 = _mid_data_in_44_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_44_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_68 = _mid_data_in_44_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_44_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_69 = _mid_data_in_44_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_44_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_70 = _mid_data_in_44_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_44_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_71 = _mid_data_in_44_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_44_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_72 = _mid_data_in_44_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_44_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_73 = _mid_data_in_44_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_44_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_74 = _mid_data_in_44_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_44_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_75 = _mid_data_in_44_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_44_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_76 = _mid_data_in_44_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_44_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_77 = _mid_data_in_44_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_44_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_78 = _mid_data_in_44_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_44_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_44_tkeep_T_79 = _mid_data_in_44_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_44_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_177 = _T_180 < 32'h10 ? _mid_data_in_44_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_178 = _T_180 < 32'h10 & _mid_data_in_44_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_44_tdata = 32'h2c >= mid_count ? _GEN_177 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_44_tkeep = 32'h2c >= mid_count & _GEN_178; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_184 = 32'h2d - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_45_tdata_T_2 = 32'h0 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_6 = 32'h1 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_10 = 32'h2 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_14 = 32'h3 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_18 = 32'h4 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_22 = 32'h5 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_26 = 32'h6 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_30 = 32'h7 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_34 = 32'h8 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_38 = 32'h9 == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_42 = 32'ha == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_46 = 32'hb == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_50 = 32'hc == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_54 = 32'hd == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_58 = 32'he == _T_184; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_45_tdata_T_62 = 32'hf == _T_184; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_45_tdata_T_64 = _mid_data_in_45_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_65 = _mid_data_in_45_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_45_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_66 = _mid_data_in_45_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_45_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_67 = _mid_data_in_45_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_45_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_68 = _mid_data_in_45_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_45_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_69 = _mid_data_in_45_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_45_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_70 = _mid_data_in_45_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_45_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_71 = _mid_data_in_45_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_45_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_72 = _mid_data_in_45_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_45_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_73 = _mid_data_in_45_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_45_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_74 = _mid_data_in_45_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_45_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_75 = _mid_data_in_45_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_45_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_76 = _mid_data_in_45_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_45_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_77 = _mid_data_in_45_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_45_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_78 = _mid_data_in_45_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_45_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_45_tdata_T_79 = _mid_data_in_45_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_45_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_65 = _mid_data_in_45_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_45_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_66 = _mid_data_in_45_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_45_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_67 = _mid_data_in_45_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_45_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_68 = _mid_data_in_45_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_45_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_69 = _mid_data_in_45_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_45_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_70 = _mid_data_in_45_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_45_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_71 = _mid_data_in_45_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_45_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_72 = _mid_data_in_45_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_45_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_73 = _mid_data_in_45_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_45_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_74 = _mid_data_in_45_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_45_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_75 = _mid_data_in_45_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_45_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_76 = _mid_data_in_45_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_45_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_77 = _mid_data_in_45_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_45_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_78 = _mid_data_in_45_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_45_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_45_tkeep_T_79 = _mid_data_in_45_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_45_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_181 = _T_184 < 32'h10 ? _mid_data_in_45_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_182 = _T_184 < 32'h10 & _mid_data_in_45_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_45_tdata = 32'h2d >= mid_count ? _GEN_181 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_45_tkeep = 32'h2d >= mid_count & _GEN_182; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_188 = 32'h2e - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_46_tdata_T_2 = 32'h0 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_6 = 32'h1 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_10 = 32'h2 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_14 = 32'h3 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_18 = 32'h4 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_22 = 32'h5 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_26 = 32'h6 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_30 = 32'h7 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_34 = 32'h8 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_38 = 32'h9 == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_42 = 32'ha == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_46 = 32'hb == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_50 = 32'hc == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_54 = 32'hd == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_58 = 32'he == _T_188; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_46_tdata_T_62 = 32'hf == _T_188; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_46_tdata_T_64 = _mid_data_in_46_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_65 = _mid_data_in_46_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_46_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_66 = _mid_data_in_46_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_46_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_67 = _mid_data_in_46_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_46_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_68 = _mid_data_in_46_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_46_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_69 = _mid_data_in_46_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_46_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_70 = _mid_data_in_46_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_46_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_71 = _mid_data_in_46_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_46_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_72 = _mid_data_in_46_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_46_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_73 = _mid_data_in_46_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_46_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_74 = _mid_data_in_46_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_46_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_75 = _mid_data_in_46_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_46_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_76 = _mid_data_in_46_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_46_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_77 = _mid_data_in_46_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_46_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_78 = _mid_data_in_46_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_46_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_46_tdata_T_79 = _mid_data_in_46_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_46_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_65 = _mid_data_in_46_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_46_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_66 = _mid_data_in_46_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_46_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_67 = _mid_data_in_46_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_46_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_68 = _mid_data_in_46_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_46_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_69 = _mid_data_in_46_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_46_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_70 = _mid_data_in_46_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_46_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_71 = _mid_data_in_46_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_46_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_72 = _mid_data_in_46_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_46_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_73 = _mid_data_in_46_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_46_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_74 = _mid_data_in_46_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_46_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_75 = _mid_data_in_46_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_46_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_76 = _mid_data_in_46_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_46_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_77 = _mid_data_in_46_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_46_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_78 = _mid_data_in_46_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_46_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_46_tkeep_T_79 = _mid_data_in_46_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_46_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_185 = _T_188 < 32'h10 ? _mid_data_in_46_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_186 = _T_188 < 32'h10 & _mid_data_in_46_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_46_tdata = 32'h2e >= mid_count ? _GEN_185 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_46_tkeep = 32'h2e >= mid_count & _GEN_186; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [31:0] _T_192 = 32'h2f - mid_count; // @[bfs_remote.scala 71:19]
  wire  _mid_data_in_47_tdata_T_2 = 32'h0 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_6 = 32'h1 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_10 = 32'h2 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_14 = 32'h3 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_18 = 32'h4 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_22 = 32'h5 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_26 = 32'h6 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_30 = 32'h7 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_34 = 32'h8 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_38 = 32'h9 == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_42 = 32'ha == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_46 = 32'hb == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_50 = 32'hc == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_54 = 32'hd == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_58 = 32'he == _T_192; // @[bfs_remote.scala 73:23]
  wire  _mid_data_in_47_tdata_T_62 = 32'hf == _T_192; // @[bfs_remote.scala 73:23]
  wire [31:0] _mid_data_in_47_tdata_T_64 = _mid_data_in_47_tdata_T_62 ? sorted_in_m_axis_tdata[511:480] : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_65 = _mid_data_in_47_tdata_T_58 ? sorted_in_m_axis_tdata[479:448] :
    _mid_data_in_47_tdata_T_64; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_66 = _mid_data_in_47_tdata_T_54 ? sorted_in_m_axis_tdata[447:416] :
    _mid_data_in_47_tdata_T_65; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_67 = _mid_data_in_47_tdata_T_50 ? sorted_in_m_axis_tdata[415:384] :
    _mid_data_in_47_tdata_T_66; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_68 = _mid_data_in_47_tdata_T_46 ? sorted_in_m_axis_tdata[383:352] :
    _mid_data_in_47_tdata_T_67; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_69 = _mid_data_in_47_tdata_T_42 ? sorted_in_m_axis_tdata[351:320] :
    _mid_data_in_47_tdata_T_68; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_70 = _mid_data_in_47_tdata_T_38 ? sorted_in_m_axis_tdata[319:288] :
    _mid_data_in_47_tdata_T_69; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_71 = _mid_data_in_47_tdata_T_34 ? sorted_in_m_axis_tdata[287:256] :
    _mid_data_in_47_tdata_T_70; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_72 = _mid_data_in_47_tdata_T_30 ? sorted_in_m_axis_tdata[255:224] :
    _mid_data_in_47_tdata_T_71; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_73 = _mid_data_in_47_tdata_T_26 ? sorted_in_m_axis_tdata[223:192] :
    _mid_data_in_47_tdata_T_72; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_74 = _mid_data_in_47_tdata_T_22 ? sorted_in_m_axis_tdata[191:160] :
    _mid_data_in_47_tdata_T_73; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_75 = _mid_data_in_47_tdata_T_18 ? sorted_in_m_axis_tdata[159:128] :
    _mid_data_in_47_tdata_T_74; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_76 = _mid_data_in_47_tdata_T_14 ? sorted_in_m_axis_tdata[127:96] :
    _mid_data_in_47_tdata_T_75; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_77 = _mid_data_in_47_tdata_T_10 ? sorted_in_m_axis_tdata[95:64] :
    _mid_data_in_47_tdata_T_76; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_78 = _mid_data_in_47_tdata_T_6 ? sorted_in_m_axis_tdata[63:32] :
    _mid_data_in_47_tdata_T_77; // @[Mux.scala 98:16]
  wire [31:0] _mid_data_in_47_tdata_T_79 = _mid_data_in_47_tdata_T_2 ? sorted_in_m_axis_tdata[31:0] :
    _mid_data_in_47_tdata_T_78; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_65 = _mid_data_in_47_tdata_T_58 ? sorted_in_m_axis_tkeep[14] :
    _mid_data_in_47_tdata_T_62 & sorted_in_m_axis_tkeep[15]; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_66 = _mid_data_in_47_tdata_T_54 ? sorted_in_m_axis_tkeep[13] :
    _mid_data_in_47_tkeep_T_65; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_67 = _mid_data_in_47_tdata_T_50 ? sorted_in_m_axis_tkeep[12] :
    _mid_data_in_47_tkeep_T_66; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_68 = _mid_data_in_47_tdata_T_46 ? sorted_in_m_axis_tkeep[11] :
    _mid_data_in_47_tkeep_T_67; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_69 = _mid_data_in_47_tdata_T_42 ? sorted_in_m_axis_tkeep[10] :
    _mid_data_in_47_tkeep_T_68; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_70 = _mid_data_in_47_tdata_T_38 ? sorted_in_m_axis_tkeep[9] : _mid_data_in_47_tkeep_T_69
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_71 = _mid_data_in_47_tdata_T_34 ? sorted_in_m_axis_tkeep[8] : _mid_data_in_47_tkeep_T_70
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_72 = _mid_data_in_47_tdata_T_30 ? sorted_in_m_axis_tkeep[7] : _mid_data_in_47_tkeep_T_71
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_73 = _mid_data_in_47_tdata_T_26 ? sorted_in_m_axis_tkeep[6] : _mid_data_in_47_tkeep_T_72
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_74 = _mid_data_in_47_tdata_T_22 ? sorted_in_m_axis_tkeep[5] : _mid_data_in_47_tkeep_T_73
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_75 = _mid_data_in_47_tdata_T_18 ? sorted_in_m_axis_tkeep[4] : _mid_data_in_47_tkeep_T_74
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_76 = _mid_data_in_47_tdata_T_14 ? sorted_in_m_axis_tkeep[3] : _mid_data_in_47_tkeep_T_75
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_77 = _mid_data_in_47_tdata_T_10 ? sorted_in_m_axis_tkeep[2] : _mid_data_in_47_tkeep_T_76
    ; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_78 = _mid_data_in_47_tdata_T_6 ? sorted_in_m_axis_tkeep[1] : _mid_data_in_47_tkeep_T_77; // @[Mux.scala 98:16]
  wire  _mid_data_in_47_tkeep_T_79 = _mid_data_in_47_tdata_T_2 ? sorted_in_m_axis_tkeep[0] : _mid_data_in_47_tkeep_T_78; // @[Mux.scala 98:16]
  wire [31:0] _GEN_189 = _T_192 < 32'h10 ? _mid_data_in_47_tdata_T_79 : 32'h0; // @[bfs_remote.scala 71:39 bfs_remote.scala 72:19 bfs_remote.scala 79:19]
  wire  _GEN_190 = _T_192 < 32'h10 & _mid_data_in_47_tkeep_T_79; // @[bfs_remote.scala 71:39 bfs_remote.scala 75:19 bfs_remote.scala 80:19]
  wire [31:0] mid_data_in_47_tdata = 32'h2f >= mid_count ? _GEN_189 : 32'h0; // @[bfs_remote.scala 70:29 bfs_remote.scala 67:17]
  wire  mid_data_in_47_tkeep = 32'h2f >= mid_count & _GEN_190; // @[bfs_remote.scala 70:29 bfs_remote.scala 68:17]
  wire [63:0] _io_out_bits_tkeep_T = out_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire  _T_194 = mid_m_axis_tvalid; // @[bfs_remote.scala 95:35]
  wire  _T_195 = mid_count >= 32'h10; // @[bfs_remote.scala 96:21]
  wire  _T_196 = _T_195 | io_flush; // @[bfs_remote.scala 97:5]
  wire [15:0] _GEN_194 = _T_195 | io_flush ? mid_m_axis_tkeep[15:0] : 16'h0; // @[bfs_remote.scala 97:17 bfs_remote.scala 99:27 bfs_remote.scala 93:23]
  wire [511:0] _GEN_195 = _T_195 | io_flush ? mid_m_axis_tdata[511:0] : 512'h0; // @[bfs_remote.scala 97:17 bfs_remote.scala 100:27 bfs_remote.scala 94:23]
  wire [15:0] _GEN_197 = mid_m_axis_tvalid ? _GEN_194 : 16'h0; // @[bfs_remote.scala 95:38 bfs_remote.scala 93:23]
  wire  _mid_io_m_axis_tready_T = out_s_axis_tready & out_s_axis_tvalid; // @[bfs_remote.scala 106:49]
  wire  _mid_io_m_axis_tready_T_1 = mid_count < 32'h10; // @[bfs_remote.scala 106:110]
  wire  _mid_io_s_axis_tvalid_T = sorted_in_m_axis_tvalid; // @[bfs_remote.scala 107:60]
  wire  _mid_io_s_axis_tvalid_T_3 = _mid_io_m_axis_tready_T & mid_count > 32'h10; // @[bfs_remote.scala 108:50]
  wire  _T_199 = out_s_axis_tvalid; // @[bfs_remote.scala 113:39]
  wire [255:0] mid_io_s_axis_tdata_lo_lo = {mid_data_in_23_tdata,mid_data_in_22_tdata,mid_data_in_21_tdata,
    mid_data_in_20_tdata,mid_data_in_19_tdata,mid_data_in_18_tdata,mid_data_in_17_tdata,mid_data_in_16_tdata}; // @[bfs_remote.scala 118:96]
  wire [511:0] mid_io_s_axis_tdata_lo = {mid_data_in_31_tdata,mid_data_in_30_tdata,mid_data_in_29_tdata,
    mid_data_in_28_tdata,mid_data_in_27_tdata,mid_data_in_26_tdata,mid_data_in_25_tdata,mid_data_in_24_tdata,
    mid_io_s_axis_tdata_lo_lo}; // @[bfs_remote.scala 118:96]
  wire [255:0] mid_io_s_axis_tdata_hi_lo = {mid_data_in_39_tdata,mid_data_in_38_tdata,mid_data_in_37_tdata,
    mid_data_in_36_tdata,mid_data_in_35_tdata,mid_data_in_34_tdata,mid_data_in_33_tdata,mid_data_in_32_tdata}; // @[bfs_remote.scala 118:96]
  wire [1023:0] _mid_io_s_axis_tdata_T = {mid_data_in_47_tdata,mid_data_in_46_tdata,mid_data_in_45_tdata,
    mid_data_in_44_tdata,mid_data_in_43_tdata,mid_data_in_42_tdata,mid_data_in_41_tdata,mid_data_in_40_tdata,
    mid_io_s_axis_tdata_hi_lo,mid_io_s_axis_tdata_lo}; // @[bfs_remote.scala 118:96]
  wire [7:0] mid_io_s_axis_tkeep_lo_lo = {mid_data_in_23_tkeep,mid_data_in_22_tkeep,mid_data_in_21_tkeep,
    mid_data_in_20_tkeep,mid_data_in_19_tkeep,mid_data_in_18_tkeep,mid_data_in_17_tkeep,mid_data_in_16_tkeep}; // @[bfs_remote.scala 119:96]
  wire [15:0] mid_io_s_axis_tkeep_lo = {mid_data_in_31_tkeep,mid_data_in_30_tkeep,mid_data_in_29_tkeep,
    mid_data_in_28_tkeep,mid_data_in_27_tkeep,mid_data_in_26_tkeep,mid_data_in_25_tkeep,mid_data_in_24_tkeep,
    mid_io_s_axis_tkeep_lo_lo}; // @[bfs_remote.scala 119:96]
  wire [7:0] mid_io_s_axis_tkeep_hi_lo = {mid_data_in_39_tkeep,mid_data_in_38_tkeep,mid_data_in_37_tkeep,
    mid_data_in_36_tkeep,mid_data_in_35_tkeep,mid_data_in_34_tkeep,mid_data_in_33_tkeep,mid_data_in_32_tkeep}; // @[bfs_remote.scala 119:96]
  wire [31:0] _mid_io_s_axis_tkeep_T = {mid_data_in_47_tkeep,mid_data_in_46_tkeep,mid_data_in_45_tkeep,
    mid_data_in_44_tkeep,mid_data_in_43_tkeep,mid_data_in_42_tkeep,mid_data_in_41_tkeep,mid_data_in_40_tkeep,
    mid_io_s_axis_tkeep_hi_lo,mid_io_s_axis_tkeep_lo}; // @[bfs_remote.scala 119:96]
  wire [1023:0] _GEN_199 = _mid_io_m_axis_tready_T_1 ? {{512'd0}, sorted_in_m_axis_tdata} : _mid_io_s_axis_tdata_T; // @[bfs_remote.scala 114:31 bfs_remote.scala 115:31 bfs_remote.scala 118:31]
  wire [63:0] _GEN_200 = _mid_io_m_axis_tready_T_1 ? sorted_in_m_axis_tkeep : {{32'd0}, _mid_io_s_axis_tkeep_T}; // @[bfs_remote.scala 114:31 bfs_remote.scala 116:31 bfs_remote.scala 119:31]
  wire [191:0] mid_io_s_axis_tdata_lo_lo_lo_1 = {mid_data_in_5_tdata,mid_data_in_4_tdata,mid_data_in_3_tdata,
    mid_data_in_2_tdata,mid_data_in_1_tdata,mid_data_in_0_tdata}; // @[bfs_remote.scala 122:75]
  wire [383:0] mid_io_s_axis_tdata_lo_lo_1 = {mid_data_in_11_tdata,mid_data_in_10_tdata,mid_data_in_9_tdata,
    mid_data_in_8_tdata,mid_data_in_7_tdata,mid_data_in_6_tdata,mid_io_s_axis_tdata_lo_lo_lo_1}; // @[bfs_remote.scala 122:75]
  wire [191:0] mid_io_s_axis_tdata_lo_hi_lo_1 = {mid_data_in_17_tdata,mid_data_in_16_tdata,mid_data_in_15_tdata,
    mid_data_in_14_tdata,mid_data_in_13_tdata,mid_data_in_12_tdata}; // @[bfs_remote.scala 122:75]
  wire [767:0] mid_io_s_axis_tdata_lo_1 = {mid_data_in_23_tdata,mid_data_in_22_tdata,mid_data_in_21_tdata,
    mid_data_in_20_tdata,mid_data_in_19_tdata,mid_data_in_18_tdata,mid_io_s_axis_tdata_lo_hi_lo_1,
    mid_io_s_axis_tdata_lo_lo_1}; // @[bfs_remote.scala 122:75]
  wire [191:0] mid_io_s_axis_tdata_hi_lo_lo_1 = {mid_data_in_29_tdata,mid_data_in_28_tdata,mid_data_in_27_tdata,
    mid_data_in_26_tdata,mid_data_in_25_tdata,mid_data_in_24_tdata}; // @[bfs_remote.scala 122:75]
  wire [383:0] mid_io_s_axis_tdata_hi_lo_1 = {mid_data_in_35_tdata,mid_data_in_34_tdata,mid_data_in_33_tdata,
    mid_data_in_32_tdata,mid_data_in_31_tdata,mid_data_in_30_tdata,mid_io_s_axis_tdata_hi_lo_lo_1}; // @[bfs_remote.scala 122:75]
  wire [191:0] mid_io_s_axis_tdata_hi_hi_lo_1 = {mid_data_in_41_tdata,mid_data_in_40_tdata,mid_data_in_39_tdata,
    mid_data_in_38_tdata,mid_data_in_37_tdata,mid_data_in_36_tdata}; // @[bfs_remote.scala 122:75]
  wire [1535:0] _mid_io_s_axis_tdata_T_1 = {mid_data_in_47_tdata,mid_data_in_46_tdata,mid_data_in_45_tdata,
    mid_data_in_44_tdata,mid_data_in_43_tdata,mid_data_in_42_tdata,mid_io_s_axis_tdata_hi_hi_lo_1,
    mid_io_s_axis_tdata_hi_lo_1,mid_io_s_axis_tdata_lo_1}; // @[bfs_remote.scala 122:75]
  wire [5:0] mid_io_s_axis_tkeep_lo_lo_lo_1 = {mid_data_in_5_tkeep,mid_data_in_4_tkeep,mid_data_in_3_tkeep,
    mid_data_in_2_tkeep,mid_data_in_1_tkeep,mid_data_in_0_tkeep}; // @[bfs_remote.scala 123:75]
  wire [11:0] mid_io_s_axis_tkeep_lo_lo_1 = {mid_data_in_11_tkeep,mid_data_in_10_tkeep,mid_data_in_9_tkeep,
    mid_data_in_8_tkeep,mid_data_in_7_tkeep,mid_data_in_6_tkeep,mid_io_s_axis_tkeep_lo_lo_lo_1}; // @[bfs_remote.scala 123:75]
  wire [5:0] mid_io_s_axis_tkeep_lo_hi_lo_1 = {mid_data_in_17_tkeep,mid_data_in_16_tkeep,mid_data_in_15_tkeep,
    mid_data_in_14_tkeep,mid_data_in_13_tkeep,mid_data_in_12_tkeep}; // @[bfs_remote.scala 123:75]
  wire [23:0] mid_io_s_axis_tkeep_lo_1 = {mid_data_in_23_tkeep,mid_data_in_22_tkeep,mid_data_in_21_tkeep,
    mid_data_in_20_tkeep,mid_data_in_19_tkeep,mid_data_in_18_tkeep,mid_io_s_axis_tkeep_lo_hi_lo_1,
    mid_io_s_axis_tkeep_lo_lo_1}; // @[bfs_remote.scala 123:75]
  wire [5:0] mid_io_s_axis_tkeep_hi_lo_lo_1 = {mid_data_in_29_tkeep,mid_data_in_28_tkeep,mid_data_in_27_tkeep,
    mid_data_in_26_tkeep,mid_data_in_25_tkeep,mid_data_in_24_tkeep}; // @[bfs_remote.scala 123:75]
  wire [11:0] mid_io_s_axis_tkeep_hi_lo_1 = {mid_data_in_35_tkeep,mid_data_in_34_tkeep,mid_data_in_33_tkeep,
    mid_data_in_32_tkeep,mid_data_in_31_tkeep,mid_data_in_30_tkeep,mid_io_s_axis_tkeep_hi_lo_lo_1}; // @[bfs_remote.scala 123:75]
  wire [5:0] mid_io_s_axis_tkeep_hi_hi_lo_1 = {mid_data_in_41_tkeep,mid_data_in_40_tkeep,mid_data_in_39_tkeep,
    mid_data_in_38_tkeep,mid_data_in_37_tkeep,mid_data_in_36_tkeep}; // @[bfs_remote.scala 123:75]
  wire [47:0] _mid_io_s_axis_tkeep_T_1 = {mid_data_in_47_tkeep,mid_data_in_46_tkeep,mid_data_in_45_tkeep,
    mid_data_in_44_tkeep,mid_data_in_43_tkeep,mid_data_in_42_tkeep,mid_io_s_axis_tkeep_hi_hi_lo_1,
    mid_io_s_axis_tkeep_hi_lo_1,mid_io_s_axis_tkeep_lo_1}; // @[bfs_remote.scala 123:75]
  wire [1535:0] _GEN_201 = out_s_axis_tvalid ? {{512'd0}, _GEN_199} : _mid_io_s_axis_tdata_T_1; // @[bfs_remote.scala 113:42 bfs_remote.scala 122:29]
  wire [63:0] _GEN_202 = out_s_axis_tvalid ? _GEN_200 : {{16'd0}, _mid_io_s_axis_tkeep_T_1}; // @[bfs_remote.scala 113:42 bfs_remote.scala 123:29]
  wire [1535:0] _GEN_203 = _T_194 ? _GEN_201 : {{1024'd0}, sorted_in_m_axis_tdata}; // @[bfs_remote.scala 112:40 bfs_remote.scala 126:27]
  wire [63:0] _GEN_204 = _T_194 ? _GEN_202 : sorted_in_m_axis_tkeep; // @[bfs_remote.scala 112:40 bfs_remote.scala 127:27]
  wire [1535:0] _GEN_205 = mid_s_axis_tvalid ? _GEN_203 : 1536'h0; // @[bfs_remote.scala 111:38 bfs_remote.scala 109:23]
  wire [63:0] _GEN_206 = mid_s_axis_tvalid ? _GEN_204 : 64'h0; // @[bfs_remote.scala 111:38 bfs_remote.scala 110:23]
  wire  _T_203 = _mid_io_s_axis_tvalid_T & sorted_in_m_axis_tready; // @[bfs_remote.scala 130:44]
  wire  _T_205 = _mid_io_s_axis_tvalid_T & sorted_in_m_axis_tready & _T_199; // @[bfs_remote.scala 130:83]
  wire  _T_206 = out_s_axis_tready; // @[bfs_remote.scala 131:65]
  wire [31:0] _mid_count_T_1 = mid_count + in_count_reg; // @[bfs_remote.scala 135:30]
  wire [31:0] _mid_count_T_3 = _mid_count_T_1 - 32'h10; // @[bfs_remote.scala 135:45]
  wire [31:0] _mid_count_T_5 = mid_count - 32'h10; // @[bfs_remote.scala 141:30]
  collector_reg in ( // @[bfs_remote.scala 19:18]
    .aclk(in_aclk),
    .aresetn(in_aresetn),
    .s_axis_tdata(in_s_axis_tdata),
    .s_axis_tvalid(in_s_axis_tvalid),
    .s_axis_tkeep(in_s_axis_tkeep),
    .s_axis_tready(in_s_axis_tready),
    .s_axis_tlast(in_s_axis_tlast),
    .m_axis_tdata(in_m_axis_tdata),
    .m_axis_tvalid(in_m_axis_tvalid),
    .m_axis_tkeep(in_m_axis_tkeep),
    .m_axis_tready(in_m_axis_tready),
    .m_axis_tlast(in_m_axis_tlast)
  );
  collector_reg sorted_in ( // @[bfs_remote.scala 43:25]
    .aclk(sorted_in_aclk),
    .aresetn(sorted_in_aresetn),
    .s_axis_tdata(sorted_in_s_axis_tdata),
    .s_axis_tvalid(sorted_in_s_axis_tvalid),
    .s_axis_tkeep(sorted_in_s_axis_tkeep),
    .s_axis_tready(sorted_in_s_axis_tready),
    .s_axis_tlast(sorted_in_s_axis_tlast),
    .m_axis_tdata(sorted_in_m_axis_tdata),
    .m_axis_tvalid(sorted_in_m_axis_tvalid),
    .m_axis_tkeep(sorted_in_m_axis_tkeep),
    .m_axis_tready(sorted_in_m_axis_tready),
    .m_axis_tlast(sorted_in_m_axis_tlast)
  );
  collector_mid_reg mid ( // @[bfs_remote.scala 55:19]
    .aclk(mid_aclk),
    .aresetn(mid_aresetn),
    .s_axis_tdata(mid_s_axis_tdata),
    .s_axis_tvalid(mid_s_axis_tvalid),
    .s_axis_tkeep(mid_s_axis_tkeep),
    .s_axis_tready(mid_s_axis_tready),
    .s_axis_tlast(mid_s_axis_tlast),
    .m_axis_tdata(mid_m_axis_tdata),
    .m_axis_tvalid(mid_m_axis_tvalid),
    .m_axis_tkeep(mid_m_axis_tkeep),
    .m_axis_tready(mid_m_axis_tready),
    .m_axis_tlast(mid_m_axis_tlast)
  );
  collector_reg out ( // @[bfs_remote.scala 86:19]
    .aclk(out_aclk),
    .aresetn(out_aresetn),
    .s_axis_tdata(out_s_axis_tdata),
    .s_axis_tvalid(out_s_axis_tvalid),
    .s_axis_tkeep(out_s_axis_tkeep),
    .s_axis_tready(out_s_axis_tready),
    .s_axis_tlast(out_s_axis_tlast),
    .m_axis_tdata(out_m_axis_tdata),
    .m_axis_tvalid(out_m_axis_tvalid),
    .m_axis_tkeep(out_m_axis_tkeep),
    .m_axis_tready(out_m_axis_tready),
    .m_axis_tlast(out_m_axis_tlast)
  );
  assign io_in_ready = in_s_axis_tready; // @[bfs_remote.scala 24:15]
  assign io_out_valid = out_m_axis_tvalid; // @[bfs_remote.scala 91:16]
  assign io_out_bits_tdata = out_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_out_bits_tkeep = _io_out_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_out_bits_tlast = out_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_empty = ~(in_m_axis_tvalid | mid_m_axis_tvalid | out_m_axis_tvalid | sorted_in_m_axis_tvalid); // @[bfs_remote.scala 148:112]
  assign in_aclk = clock; // @[bfs_remote.scala 20:29]
  assign in_aresetn = ~reset; // @[bfs_remote.scala 21:20]
  assign in_s_axis_tdata = io_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign in_s_axis_tvalid = io_in_valid; // @[bfs_remote.scala 22:23]
  assign in_s_axis_tkeep = {{48'd0}, io_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign in_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign in_m_axis_tready = sorted_in_s_axis_tready | in_count_15 == 8'h0; // @[bfs_remote.scala 49:53]
  assign sorted_in_aclk = clock; // @[bfs_remote.scala 44:36]
  assign sorted_in_aresetn = ~reset; // @[bfs_remote.scala 45:27]
  assign sorted_in_s_axis_tdata = {sorted_in_io_s_axis_tdata_hi,sorted_in_io_s_axis_tdata_lo}; // @[bfs_remote.scala 48:71]
  assign sorted_in_s_axis_tvalid = in_m_axis_tvalid & in_count_15 > 8'h0; // @[bfs_remote.scala 46:53]
  assign sorted_in_s_axis_tkeep = {{48'd0}, _sorted_in_io_s_axis_tkeep_T}; // @[bfs_remote.scala 47:71]
  assign sorted_in_s_axis_tlast = 1'h0;
  assign sorted_in_m_axis_tready = mid_s_axis_tready; // @[bfs_remote.scala 147:30]
  assign mid_aclk = clock; // @[bfs_remote.scala 56:30]
  assign mid_aresetn = ~reset; // @[bfs_remote.scala 57:21]
  assign mid_s_axis_tdata = _GEN_205[1023:0];
  assign mid_s_axis_tvalid = sorted_in_m_axis_tvalid | _mid_io_s_axis_tvalid_T_3; // @[bfs_remote.scala 107:63]
  assign mid_s_axis_tkeep = {{64'd0}, _GEN_206}; // @[bfs_remote.scala 111:38 bfs_remote.scala 110:23]
  assign mid_s_axis_tlast = 1'h0;
  assign mid_m_axis_tready = out_s_axis_tready & out_s_axis_tvalid | mid_s_axis_tvalid & mid_count < 32'h10; // @[bfs_remote.scala 106:73]
  assign out_aclk = clock; // @[bfs_remote.scala 87:30]
  assign out_aresetn = ~reset; // @[bfs_remote.scala 88:21]
  assign out_s_axis_tdata = mid_m_axis_tvalid ? _GEN_195 : 512'h0; // @[bfs_remote.scala 95:38 bfs_remote.scala 94:23]
  assign out_s_axis_tvalid = mid_m_axis_tvalid & _T_196; // @[bfs_remote.scala 95:38 bfs_remote.scala 92:24]
  assign out_s_axis_tkeep = {{48'd0}, _GEN_197}; // @[bfs_remote.scala 95:38 bfs_remote.scala 93:23]
  assign out_s_axis_tlast = 1'h1; // @[bfs_remote.scala 103:23]
  assign out_m_axis_tready = io_out_ready; // @[bfs_remote.scala 89:24]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 50:29]
      in_count_reg <= 32'h0; // @[bfs_remote.scala 50:29]
    end else if (sorted_in_s_axis_tvalid & sorted_in_s_axis_tready) begin // @[bfs_remote.scala 51:75]
      in_count_reg <= {{24'd0}, in_count_15}; // @[bfs_remote.scala 52:18]
    end
    if (reset) begin // @[bfs_remote.scala 58:26]
      mid_count <= 32'h0; // @[bfs_remote.scala 58:26]
    end else if (_T_205 & out_s_axis_tready) begin // @[bfs_remote.scala 131:68]
      if (_mid_io_m_axis_tready_T_1) begin // @[bfs_remote.scala 132:27]
        mid_count <= in_count_reg; // @[bfs_remote.scala 133:17]
      end else begin
        mid_count <= _mid_count_T_3; // @[bfs_remote.scala 135:17]
      end
    end else if (_T_199 & _T_206) begin // @[bfs_remote.scala 137:77]
      if (_mid_io_m_axis_tready_T_1) begin // @[bfs_remote.scala 138:27]
        mid_count <= 32'h0; // @[bfs_remote.scala 139:17]
      end else begin
        mid_count <= _mid_count_T_5; // @[bfs_remote.scala 141:17]
      end
    end else if (_T_203) begin // @[bfs_remote.scala 143:89]
      mid_count <= _mid_count_T_1; // @[bfs_remote.scala 144:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_count_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mid_count = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [511:0] io_in_0_bits_tdata,
  input  [63:0]  io_in_0_bits_tkeep,
  input          io_in_0_bits_tlast,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [511:0] io_in_1_bits_tdata,
  input  [63:0]  io_in_1_bits_tkeep,
  input          io_in_1_bits_tlast,
  input          io_out_ready,
  output         io_out_valid,
  output [511:0] io_out_bits_tdata,
  output [63:0]  io_out_bits_tkeep,
  output         io_out_bits_tlast
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_tdata = io_in_0_valid ? io_in_0_bits_tdata : io_in_1_bits_tdata; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_tkeep = io_in_0_valid ? io_in_0_bits_tkeep : io_in_1_bits_tkeep; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_tlast = io_in_0_valid ? io_in_0_bits_tlast : io_in_1_bits_tlast; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
endmodule
module Remote_xbar(
  input          clock,
  input          reset,
  output         io_ddr_in_0_ready,
  input          io_ddr_in_0_valid,
  input  [127:0] io_ddr_in_0_bits_tdata,
  input  [3:0]   io_ddr_in_0_bits_tkeep,
  input          io_ddr_in_0_bits_tlast,
  output         io_ddr_in_1_ready,
  input          io_ddr_in_1_valid,
  input  [127:0] io_ddr_in_1_bits_tdata,
  input  [3:0]   io_ddr_in_1_bits_tkeep,
  input          io_ddr_in_1_bits_tlast,
  output         io_ddr_in_2_ready,
  input          io_ddr_in_2_valid,
  input  [127:0] io_ddr_in_2_bits_tdata,
  input  [3:0]   io_ddr_in_2_bits_tkeep,
  input          io_ddr_in_2_bits_tlast,
  output         io_ddr_in_3_ready,
  input          io_ddr_in_3_valid,
  input  [127:0] io_ddr_in_3_bits_tdata,
  input  [3:0]   io_ddr_in_3_bits_tkeep,
  input          io_ddr_in_3_bits_tlast,
  input          io_pe_out_0_ready,
  output         io_pe_out_0_valid,
  output [511:0] io_pe_out_0_bits_tdata,
  output [15:0]  io_pe_out_0_bits_tkeep,
  output         io_pe_out_0_bits_tlast,
  input          io_pe_out_1_ready,
  output         io_pe_out_1_valid,
  output [511:0] io_pe_out_1_bits_tdata,
  output [15:0]  io_pe_out_1_bits_tkeep,
  output         io_pe_out_1_bits_tlast,
  input          io_pe_out_2_ready,
  output         io_pe_out_2_valid,
  output [511:0] io_pe_out_2_bits_tdata,
  output [15:0]  io_pe_out_2_bits_tkeep,
  output         io_pe_out_2_bits_tlast,
  input          io_pe_out_3_ready,
  output         io_pe_out_3_valid,
  output [511:0] io_pe_out_3_bits_tdata,
  output [15:0]  io_pe_out_3_bits_tkeep,
  output         io_pe_out_3_bits_tlast,
  input          io_pe_out_4_ready,
  output         io_pe_out_4_valid,
  output [511:0] io_pe_out_4_bits_tdata,
  output [15:0]  io_pe_out_4_bits_tkeep,
  output         io_pe_out_4_bits_tlast,
  input          io_pe_out_5_ready,
  output         io_pe_out_5_valid,
  output [511:0] io_pe_out_5_bits_tdata,
  output [15:0]  io_pe_out_5_bits_tkeep,
  output         io_pe_out_5_bits_tlast,
  input          io_pe_out_6_ready,
  output         io_pe_out_6_valid,
  output [511:0] io_pe_out_6_bits_tdata,
  output [15:0]  io_pe_out_6_bits_tkeep,
  output         io_pe_out_6_bits_tlast,
  input          io_pe_out_7_ready,
  output         io_pe_out_7_valid,
  output [511:0] io_pe_out_7_bits_tdata,
  output [15:0]  io_pe_out_7_bits_tkeep,
  output         io_pe_out_7_bits_tlast,
  input          io_pe_out_8_ready,
  output         io_pe_out_8_valid,
  output [511:0] io_pe_out_8_bits_tdata,
  output [15:0]  io_pe_out_8_bits_tkeep,
  output         io_pe_out_8_bits_tlast,
  input          io_pe_out_9_ready,
  output         io_pe_out_9_valid,
  output [511:0] io_pe_out_9_bits_tdata,
  output [15:0]  io_pe_out_9_bits_tkeep,
  output         io_pe_out_9_bits_tlast,
  input          io_pe_out_10_ready,
  output         io_pe_out_10_valid,
  output [511:0] io_pe_out_10_bits_tdata,
  output [15:0]  io_pe_out_10_bits_tkeep,
  output         io_pe_out_10_bits_tlast,
  input          io_pe_out_11_ready,
  output         io_pe_out_11_valid,
  output [511:0] io_pe_out_11_bits_tdata,
  output [15:0]  io_pe_out_11_bits_tkeep,
  output         io_pe_out_11_bits_tlast,
  input          io_pe_out_12_ready,
  output         io_pe_out_12_valid,
  output [511:0] io_pe_out_12_bits_tdata,
  output [15:0]  io_pe_out_12_bits_tkeep,
  output         io_pe_out_12_bits_tlast,
  input          io_pe_out_13_ready,
  output         io_pe_out_13_valid,
  output [511:0] io_pe_out_13_bits_tdata,
  output [15:0]  io_pe_out_13_bits_tkeep,
  output         io_pe_out_13_bits_tlast,
  input          io_pe_out_14_ready,
  output         io_pe_out_14_valid,
  output [511:0] io_pe_out_14_bits_tdata,
  output [15:0]  io_pe_out_14_bits_tkeep,
  output         io_pe_out_14_bits_tlast,
  input          io_pe_out_15_ready,
  output         io_pe_out_15_valid,
  output [511:0] io_pe_out_15_bits_tdata,
  output [15:0]  io_pe_out_15_bits_tkeep,
  output         io_pe_out_15_bits_tlast,
  input          io_remote_out_0_ready,
  output         io_remote_out_0_valid,
  output [511:0] io_remote_out_0_bits_tdata,
  output [15:0]  io_remote_out_0_bits_tkeep,
  input          io_remote_out_1_ready,
  output         io_remote_out_1_valid,
  output [511:0] io_remote_out_1_bits_tdata,
  output [15:0]  io_remote_out_1_bits_tkeep,
  input          io_remote_out_2_ready,
  output         io_remote_out_2_valid,
  output [511:0] io_remote_out_2_bits_tdata,
  output [15:0]  io_remote_out_2_bits_tkeep,
  input          io_remote_out_3_ready,
  output         io_remote_out_3_valid,
  output [511:0] io_remote_out_3_bits_tdata,
  output [15:0]  io_remote_out_3_bits_tkeep,
  output         io_remote_in_ready,
  input          io_remote_in_valid,
  input  [511:0] io_remote_in_bits_tdata,
  input  [15:0]  io_remote_in_bits_tkeep,
  input  [1:0]   io_local_fpga_id,
  input          io_flush,
  input          io_signal
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  combiner_level0_aclk; // @[bfs_remote.scala 628:31]
  wire  combiner_level0_aresetn; // @[bfs_remote.scala 628:31]
  wire [511:0] combiner_level0_s_axis_tdata; // @[bfs_remote.scala 628:31]
  wire [3:0] combiner_level0_s_axis_tvalid; // @[bfs_remote.scala 628:31]
  wire [63:0] combiner_level0_s_axis_tkeep; // @[bfs_remote.scala 628:31]
  wire [3:0] combiner_level0_s_axis_tready; // @[bfs_remote.scala 628:31]
  wire [3:0] combiner_level0_s_axis_tlast; // @[bfs_remote.scala 628:31]
  wire [3:0] combiner_level0_s_axis_tid; // @[bfs_remote.scala 628:31]
  wire [511:0] combiner_level0_m_axis_tdata; // @[bfs_remote.scala 628:31]
  wire  combiner_level0_m_axis_tvalid; // @[bfs_remote.scala 628:31]
  wire [63:0] combiner_level0_m_axis_tkeep; // @[bfs_remote.scala 628:31]
  wire  combiner_level0_m_axis_tready; // @[bfs_remote.scala 628:31]
  wire  combiner_level0_m_axis_tlast; // @[bfs_remote.scala 628:31]
  wire  combiner_level0_m_axis_tid; // @[bfs_remote.scala 628:31]
  wire  frontend_aclk; // @[bfs_remote.scala 640:24]
  wire  frontend_aresetn; // @[bfs_remote.scala 640:24]
  wire [511:0] frontend_s_axis_tdata; // @[bfs_remote.scala 640:24]
  wire  frontend_s_axis_tvalid; // @[bfs_remote.scala 640:24]
  wire [63:0] frontend_s_axis_tkeep; // @[bfs_remote.scala 640:24]
  wire  frontend_s_axis_tready; // @[bfs_remote.scala 640:24]
  wire  frontend_s_axis_tlast; // @[bfs_remote.scala 640:24]
  wire [511:0] frontend_m_axis_tdata; // @[bfs_remote.scala 640:24]
  wire  frontend_m_axis_tvalid; // @[bfs_remote.scala 640:24]
  wire [63:0] frontend_m_axis_tkeep; // @[bfs_remote.scala 640:24]
  wire  frontend_m_axis_tready; // @[bfs_remote.scala 640:24]
  wire  frontend_m_axis_tlast; // @[bfs_remote.scala 640:24]
  wire  xbar_level0_aclk; // @[bfs_remote.scala 649:27]
  wire  xbar_level0_aresetn; // @[bfs_remote.scala 649:27]
  wire [511:0] xbar_level0_s_axis_tdata; // @[bfs_remote.scala 649:27]
  wire  xbar_level0_s_axis_tvalid; // @[bfs_remote.scala 649:27]
  wire [63:0] xbar_level0_s_axis_tkeep; // @[bfs_remote.scala 649:27]
  wire  xbar_level0_s_axis_tready; // @[bfs_remote.scala 649:27]
  wire  xbar_level0_s_axis_tlast; // @[bfs_remote.scala 649:27]
  wire  xbar_level0_s_axis_tid; // @[bfs_remote.scala 649:27]
  wire [2559:0] xbar_level0_m_axis_tdata; // @[bfs_remote.scala 649:27]
  wire [4:0] xbar_level0_m_axis_tvalid; // @[bfs_remote.scala 649:27]
  wire [319:0] xbar_level0_m_axis_tkeep; // @[bfs_remote.scala 649:27]
  wire [4:0] xbar_level0_m_axis_tready; // @[bfs_remote.scala 649:27]
  wire [4:0] xbar_level0_m_axis_tlast; // @[bfs_remote.scala 649:27]
  wire [4:0] xbar_level0_m_axis_tid; // @[bfs_remote.scala 649:27]
  wire  collector_clock; // @[bfs_remote.scala 682:25]
  wire  collector_reset; // @[bfs_remote.scala 682:25]
  wire  collector_io_in_ready; // @[bfs_remote.scala 682:25]
  wire  collector_io_in_valid; // @[bfs_remote.scala 682:25]
  wire [511:0] collector_io_in_bits_tdata; // @[bfs_remote.scala 682:25]
  wire [15:0] collector_io_in_bits_tkeep; // @[bfs_remote.scala 682:25]
  wire  collector_io_out_ready; // @[bfs_remote.scala 682:25]
  wire  collector_io_out_valid; // @[bfs_remote.scala 682:25]
  wire [511:0] collector_io_out_bits_tdata; // @[bfs_remote.scala 682:25]
  wire [15:0] collector_io_out_bits_tkeep; // @[bfs_remote.scala 682:25]
  wire  collector_io_out_bits_tlast; // @[bfs_remote.scala 682:25]
  wire  collector_io_flush; // @[bfs_remote.scala 682:25]
  wire  collector_io_empty; // @[bfs_remote.scala 682:25]
  wire  buffer1_s_axis_aclk; // @[bfs_remote.scala 690:23]
  wire  buffer1_s_axis_aresetn; // @[bfs_remote.scala 690:23]
  wire [511:0] buffer1_s_axis_tdata; // @[bfs_remote.scala 690:23]
  wire  buffer1_s_axis_tvalid; // @[bfs_remote.scala 690:23]
  wire [63:0] buffer1_s_axis_tkeep; // @[bfs_remote.scala 690:23]
  wire  buffer1_s_axis_tready; // @[bfs_remote.scala 690:23]
  wire  buffer1_s_axis_tlast; // @[bfs_remote.scala 690:23]
  wire  buffer1_s_axis_tid; // @[bfs_remote.scala 690:23]
  wire [511:0] buffer1_m_axis_tdata; // @[bfs_remote.scala 690:23]
  wire  buffer1_m_axis_tvalid; // @[bfs_remote.scala 690:23]
  wire [63:0] buffer1_m_axis_tkeep; // @[bfs_remote.scala 690:23]
  wire  buffer1_m_axis_tready; // @[bfs_remote.scala 690:23]
  wire  buffer1_m_axis_tlast; // @[bfs_remote.scala 690:23]
  wire  buffer1_m_axis_tid; // @[bfs_remote.scala 690:23]
  wire  remote_in_reg_aclk; // @[bfs_remote.scala 697:29]
  wire  remote_in_reg_aresetn; // @[bfs_remote.scala 697:29]
  wire [511:0] remote_in_reg_s_axis_tdata; // @[bfs_remote.scala 697:29]
  wire  remote_in_reg_s_axis_tvalid; // @[bfs_remote.scala 697:29]
  wire [63:0] remote_in_reg_s_axis_tkeep; // @[bfs_remote.scala 697:29]
  wire  remote_in_reg_s_axis_tready; // @[bfs_remote.scala 697:29]
  wire  remote_in_reg_s_axis_tlast; // @[bfs_remote.scala 697:29]
  wire [511:0] remote_in_reg_m_axis_tdata; // @[bfs_remote.scala 697:29]
  wire  remote_in_reg_m_axis_tvalid; // @[bfs_remote.scala 697:29]
  wire [63:0] remote_in_reg_m_axis_tkeep; // @[bfs_remote.scala 697:29]
  wire  remote_in_reg_m_axis_tready; // @[bfs_remote.scala 697:29]
  wire  remote_in_reg_m_axis_tlast; // @[bfs_remote.scala 697:29]
  wire  switch_level1_io_in_0_ready; // @[bfs_remote.scala 704:29]
  wire  switch_level1_io_in_0_valid; // @[bfs_remote.scala 704:29]
  wire [511:0] switch_level1_io_in_0_bits_tdata; // @[bfs_remote.scala 704:29]
  wire [63:0] switch_level1_io_in_0_bits_tkeep; // @[bfs_remote.scala 704:29]
  wire  switch_level1_io_in_0_bits_tlast; // @[bfs_remote.scala 704:29]
  wire  switch_level1_io_in_1_ready; // @[bfs_remote.scala 704:29]
  wire  switch_level1_io_in_1_valid; // @[bfs_remote.scala 704:29]
  wire [511:0] switch_level1_io_in_1_bits_tdata; // @[bfs_remote.scala 704:29]
  wire [63:0] switch_level1_io_in_1_bits_tkeep; // @[bfs_remote.scala 704:29]
  wire  switch_level1_io_in_1_bits_tlast; // @[bfs_remote.scala 704:29]
  wire  switch_level1_io_out_ready; // @[bfs_remote.scala 704:29]
  wire  switch_level1_io_out_valid; // @[bfs_remote.scala 704:29]
  wire [511:0] switch_level1_io_out_bits_tdata; // @[bfs_remote.scala 704:29]
  wire [63:0] switch_level1_io_out_bits_tkeep; // @[bfs_remote.scala 704:29]
  wire  switch_level1_io_out_bits_tlast; // @[bfs_remote.scala 704:29]
  wire  mid_aclk; // @[bfs_remote.scala 724:19]
  wire  mid_aresetn; // @[bfs_remote.scala 724:19]
  wire [511:0] mid_s_axis_tdata; // @[bfs_remote.scala 724:19]
  wire  mid_s_axis_tvalid; // @[bfs_remote.scala 724:19]
  wire [63:0] mid_s_axis_tkeep; // @[bfs_remote.scala 724:19]
  wire  mid_s_axis_tready; // @[bfs_remote.scala 724:19]
  wire  mid_s_axis_tlast; // @[bfs_remote.scala 724:19]
  wire [511:0] mid_m_axis_tdata; // @[bfs_remote.scala 724:19]
  wire  mid_m_axis_tvalid; // @[bfs_remote.scala 724:19]
  wire [63:0] mid_m_axis_tkeep; // @[bfs_remote.scala 724:19]
  wire  mid_m_axis_tready; // @[bfs_remote.scala 724:19]
  wire  mid_m_axis_tlast; // @[bfs_remote.scala 724:19]
  wire  xbar_level1_aclk; // @[bfs_remote.scala 733:27]
  wire  xbar_level1_aresetn; // @[bfs_remote.scala 733:27]
  wire [511:0] xbar_level1_s_axis_tdata; // @[bfs_remote.scala 733:27]
  wire  xbar_level1_s_axis_tvalid; // @[bfs_remote.scala 733:27]
  wire [63:0] xbar_level1_s_axis_tkeep; // @[bfs_remote.scala 733:27]
  wire  xbar_level1_s_axis_tready; // @[bfs_remote.scala 733:27]
  wire  xbar_level1_s_axis_tlast; // @[bfs_remote.scala 733:27]
  wire  xbar_level1_s_axis_tid; // @[bfs_remote.scala 733:27]
  wire [8191:0] xbar_level1_m_axis_tdata; // @[bfs_remote.scala 733:27]
  wire [15:0] xbar_level1_m_axis_tvalid; // @[bfs_remote.scala 733:27]
  wire [1023:0] xbar_level1_m_axis_tkeep; // @[bfs_remote.scala 733:27]
  wire [15:0] xbar_level1_m_axis_tready; // @[bfs_remote.scala 733:27]
  wire [15:0] xbar_level1_m_axis_tlast; // @[bfs_remote.scala 733:27]
  wire [15:0] xbar_level1_m_axis_tid; // @[bfs_remote.scala 733:27]
  wire  backend_0_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_0_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_0_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_0_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_0_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_0_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_0_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_0_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_0_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_0_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_0_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_0_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_1_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_1_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_1_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_1_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_1_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_1_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_1_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_1_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_1_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_1_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_1_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_1_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_2_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_2_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_2_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_2_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_2_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_2_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_2_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_2_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_2_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_2_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_2_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_2_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_3_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_3_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_3_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_3_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_3_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_3_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_3_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_3_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_3_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_3_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_3_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_3_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_4_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_4_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_4_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_4_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_4_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_4_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_4_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_4_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_4_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_4_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_4_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_4_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_5_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_5_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_5_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_5_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_5_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_5_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_5_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_5_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_5_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_5_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_5_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_5_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_6_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_6_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_6_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_6_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_6_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_6_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_6_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_6_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_6_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_6_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_6_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_6_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_7_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_7_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_7_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_7_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_7_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_7_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_7_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_7_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_7_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_7_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_7_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_7_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_8_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_8_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_8_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_8_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_8_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_8_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_8_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_8_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_8_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_8_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_8_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_8_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_9_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_9_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_9_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_9_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_9_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_9_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_9_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_9_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_9_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_9_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_9_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_9_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_10_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_10_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_10_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_10_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_10_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_10_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_10_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_10_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_10_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_10_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_10_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_10_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_11_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_11_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_11_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_11_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_11_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_11_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_11_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_11_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_11_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_11_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_11_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_11_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_12_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_12_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_12_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_12_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_12_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_12_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_12_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_12_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_12_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_12_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_12_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_12_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_13_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_13_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_13_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_13_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_13_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_13_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_13_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_13_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_13_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_13_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_13_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_13_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_14_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_14_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_14_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_14_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_14_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_14_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_14_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_14_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_14_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_14_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_14_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_14_m_axis_tlast; // @[bfs_remote.scala 741:43]
  wire  backend_15_aclk; // @[bfs_remote.scala 741:43]
  wire  backend_15_aresetn; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_15_s_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_15_s_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_15_s_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_15_s_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_15_s_axis_tlast; // @[bfs_remote.scala 741:43]
  wire [511:0] backend_15_m_axis_tdata; // @[bfs_remote.scala 741:43]
  wire  backend_15_m_axis_tvalid; // @[bfs_remote.scala 741:43]
  wire [63:0] backend_15_m_axis_tkeep; // @[bfs_remote.scala 741:43]
  wire  backend_15_m_axis_tready; // @[bfs_remote.scala 741:43]
  wire  backend_15_m_axis_tlast; // @[bfs_remote.scala 741:43]
  reg [1:0] local_fpga_id; // @[bfs_remote.scala 625:30]
  wire [255:0] combiner_level0_io_s_axis_tdata_lo = {io_ddr_in_1_bits_tdata,io_ddr_in_0_bits_tdata}; // @[bfs_remote.scala 631:103]
  wire [255:0] combiner_level0_io_s_axis_tdata_hi = {io_ddr_in_3_bits_tdata,io_ddr_in_2_bits_tdata}; // @[bfs_remote.scala 631:103]
  wire  _combiner_level0_io_s_axis_tkeep_T_4 = io_ddr_in_0_bits_tkeep[0] & io_ddr_in_0_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_5 = io_ddr_in_0_bits_tkeep[1] & io_ddr_in_0_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_6 = io_ddr_in_0_bits_tkeep[2] & io_ddr_in_0_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_7 = io_ddr_in_0_bits_tkeep[3] & io_ddr_in_0_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_12 = io_ddr_in_1_bits_tkeep[0] & io_ddr_in_1_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_13 = io_ddr_in_1_bits_tkeep[1] & io_ddr_in_1_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_14 = io_ddr_in_1_bits_tkeep[2] & io_ddr_in_1_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_15 = io_ddr_in_1_bits_tkeep[3] & io_ddr_in_1_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_20 = io_ddr_in_2_bits_tkeep[0] & io_ddr_in_2_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_21 = io_ddr_in_2_bits_tkeep[1] & io_ddr_in_2_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_22 = io_ddr_in_2_bits_tkeep[2] & io_ddr_in_2_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_23 = io_ddr_in_2_bits_tkeep[3] & io_ddr_in_2_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_28 = io_ddr_in_3_bits_tkeep[0] & io_ddr_in_3_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_29 = io_ddr_in_3_bits_tkeep[1] & io_ddr_in_3_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_30 = io_ddr_in_3_bits_tkeep[2] & io_ddr_in_3_valid; // @[bfs_remote.scala 632:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_31 = io_ddr_in_3_bits_tkeep[3] & io_ddr_in_3_valid; // @[bfs_remote.scala 632:125]
  wire [7:0] combiner_level0_io_s_axis_tkeep_lo = {_combiner_level0_io_s_axis_tkeep_T_15,
    _combiner_level0_io_s_axis_tkeep_T_14,_combiner_level0_io_s_axis_tkeep_T_13,_combiner_level0_io_s_axis_tkeep_T_12,
    _combiner_level0_io_s_axis_tkeep_T_7,_combiner_level0_io_s_axis_tkeep_T_6,_combiner_level0_io_s_axis_tkeep_T_5,
    _combiner_level0_io_s_axis_tkeep_T_4}; // @[bfs_remote.scala 633:33]
  wire [15:0] _combiner_level0_io_s_axis_tkeep_T_32 = {_combiner_level0_io_s_axis_tkeep_T_31,
    _combiner_level0_io_s_axis_tkeep_T_30,_combiner_level0_io_s_axis_tkeep_T_29,_combiner_level0_io_s_axis_tkeep_T_28,
    _combiner_level0_io_s_axis_tkeep_T_23,_combiner_level0_io_s_axis_tkeep_T_22,_combiner_level0_io_s_axis_tkeep_T_21,
    _combiner_level0_io_s_axis_tkeep_T_20,combiner_level0_io_s_axis_tkeep_lo}; // @[bfs_remote.scala 633:33]
  wire [1:0] combiner_level0_io_s_axis_tlast_lo = {io_ddr_in_1_bits_tlast,io_ddr_in_0_bits_tlast}; // @[bfs_remote.scala 634:103]
  wire [1:0] combiner_level0_io_s_axis_tlast_hi = {io_ddr_in_3_bits_tlast,io_ddr_in_2_bits_tlast}; // @[bfs_remote.scala 634:103]
  wire  _combiner_level0_io_s_axis_tvalid_T_2 = io_ddr_in_0_valid | io_ddr_in_1_valid | io_ddr_in_2_valid |
    io_ddr_in_3_valid; // @[bfs_remote.scala 635:104]
  wire [1:0] combiner_level0_io_s_axis_tvalid_lo = {_combiner_level0_io_s_axis_tvalid_T_2,
    _combiner_level0_io_s_axis_tvalid_T_2}; // @[bfs_remote.scala 635:116]
  wire  _xbar_level0_io_s_axis_tkeep_T_64 = frontend_m_axis_tkeep[0] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_65 = frontend_m_axis_tkeep[1] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_66 = frontend_m_axis_tkeep[2] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_67 = frontend_m_axis_tkeep[3] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_68 = frontend_m_axis_tkeep[4] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_69 = frontend_m_axis_tkeep[5] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_70 = frontend_m_axis_tkeep[6] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_71 = frontend_m_axis_tkeep[7] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_72 = frontend_m_axis_tkeep[8] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_73 = frontend_m_axis_tkeep[9] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_74 = frontend_m_axis_tkeep[10] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_75 = frontend_m_axis_tkeep[11] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_76 = frontend_m_axis_tkeep[12] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_77 = frontend_m_axis_tkeep[13] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_78 = frontend_m_axis_tkeep[14] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_79 = frontend_m_axis_tkeep[15] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_80 = frontend_m_axis_tkeep[16] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_81 = frontend_m_axis_tkeep[17] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_82 = frontend_m_axis_tkeep[18] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_83 = frontend_m_axis_tkeep[19] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_84 = frontend_m_axis_tkeep[20] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_85 = frontend_m_axis_tkeep[21] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_86 = frontend_m_axis_tkeep[22] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_87 = frontend_m_axis_tkeep[23] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_88 = frontend_m_axis_tkeep[24] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_89 = frontend_m_axis_tkeep[25] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_90 = frontend_m_axis_tkeep[26] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_91 = frontend_m_axis_tkeep[27] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_92 = frontend_m_axis_tkeep[28] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_93 = frontend_m_axis_tkeep[29] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_94 = frontend_m_axis_tkeep[30] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_95 = frontend_m_axis_tkeep[31] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_96 = frontend_m_axis_tkeep[32] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_97 = frontend_m_axis_tkeep[33] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_98 = frontend_m_axis_tkeep[34] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_99 = frontend_m_axis_tkeep[35] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_100 = frontend_m_axis_tkeep[36] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_101 = frontend_m_axis_tkeep[37] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_102 = frontend_m_axis_tkeep[38] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_103 = frontend_m_axis_tkeep[39] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_104 = frontend_m_axis_tkeep[40] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_105 = frontend_m_axis_tkeep[41] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_106 = frontend_m_axis_tkeep[42] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_107 = frontend_m_axis_tkeep[43] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_108 = frontend_m_axis_tkeep[44] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_109 = frontend_m_axis_tkeep[45] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_110 = frontend_m_axis_tkeep[46] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_111 = frontend_m_axis_tkeep[47] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_112 = frontend_m_axis_tkeep[48] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_113 = frontend_m_axis_tkeep[49] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_114 = frontend_m_axis_tkeep[50] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_115 = frontend_m_axis_tkeep[51] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_116 = frontend_m_axis_tkeep[52] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_117 = frontend_m_axis_tkeep[53] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_118 = frontend_m_axis_tkeep[54] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_119 = frontend_m_axis_tkeep[55] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_120 = frontend_m_axis_tkeep[56] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_121 = frontend_m_axis_tkeep[57] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_122 = frontend_m_axis_tkeep[58] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_123 = frontend_m_axis_tkeep[59] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_124 = frontend_m_axis_tkeep[60] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_125 = frontend_m_axis_tkeep[61] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_126 = frontend_m_axis_tkeep[62] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire  _xbar_level0_io_s_axis_tkeep_T_127 = frontend_m_axis_tkeep[63] & frontend_m_axis_tvalid; // @[bfs_remote.scala 654:88]
  wire [7:0] xbar_level0_io_s_axis_tkeep_lo_lo_lo = {_xbar_level0_io_s_axis_tkeep_T_71,_xbar_level0_io_s_axis_tkeep_T_70
    ,_xbar_level0_io_s_axis_tkeep_T_69,_xbar_level0_io_s_axis_tkeep_T_68,_xbar_level0_io_s_axis_tkeep_T_67,
    _xbar_level0_io_s_axis_tkeep_T_66,_xbar_level0_io_s_axis_tkeep_T_65,_xbar_level0_io_s_axis_tkeep_T_64}; // @[bfs_remote.scala 654:124]
  wire [15:0] xbar_level0_io_s_axis_tkeep_lo_lo = {_xbar_level0_io_s_axis_tkeep_T_79,_xbar_level0_io_s_axis_tkeep_T_78,
    _xbar_level0_io_s_axis_tkeep_T_77,_xbar_level0_io_s_axis_tkeep_T_76,_xbar_level0_io_s_axis_tkeep_T_75,
    _xbar_level0_io_s_axis_tkeep_T_74,_xbar_level0_io_s_axis_tkeep_T_73,_xbar_level0_io_s_axis_tkeep_T_72,
    xbar_level0_io_s_axis_tkeep_lo_lo_lo}; // @[bfs_remote.scala 654:124]
  wire [7:0] xbar_level0_io_s_axis_tkeep_lo_hi_lo = {_xbar_level0_io_s_axis_tkeep_T_87,_xbar_level0_io_s_axis_tkeep_T_86
    ,_xbar_level0_io_s_axis_tkeep_T_85,_xbar_level0_io_s_axis_tkeep_T_84,_xbar_level0_io_s_axis_tkeep_T_83,
    _xbar_level0_io_s_axis_tkeep_T_82,_xbar_level0_io_s_axis_tkeep_T_81,_xbar_level0_io_s_axis_tkeep_T_80}; // @[bfs_remote.scala 654:124]
  wire [31:0] xbar_level0_io_s_axis_tkeep_lo = {_xbar_level0_io_s_axis_tkeep_T_95,_xbar_level0_io_s_axis_tkeep_T_94,
    _xbar_level0_io_s_axis_tkeep_T_93,_xbar_level0_io_s_axis_tkeep_T_92,_xbar_level0_io_s_axis_tkeep_T_91,
    _xbar_level0_io_s_axis_tkeep_T_90,_xbar_level0_io_s_axis_tkeep_T_89,_xbar_level0_io_s_axis_tkeep_T_88,
    xbar_level0_io_s_axis_tkeep_lo_hi_lo,xbar_level0_io_s_axis_tkeep_lo_lo}; // @[bfs_remote.scala 654:124]
  wire [7:0] xbar_level0_io_s_axis_tkeep_hi_lo_lo = {_xbar_level0_io_s_axis_tkeep_T_103,
    _xbar_level0_io_s_axis_tkeep_T_102,_xbar_level0_io_s_axis_tkeep_T_101,_xbar_level0_io_s_axis_tkeep_T_100,
    _xbar_level0_io_s_axis_tkeep_T_99,_xbar_level0_io_s_axis_tkeep_T_98,_xbar_level0_io_s_axis_tkeep_T_97,
    _xbar_level0_io_s_axis_tkeep_T_96}; // @[bfs_remote.scala 654:124]
  wire [15:0] xbar_level0_io_s_axis_tkeep_hi_lo = {_xbar_level0_io_s_axis_tkeep_T_111,_xbar_level0_io_s_axis_tkeep_T_110
    ,_xbar_level0_io_s_axis_tkeep_T_109,_xbar_level0_io_s_axis_tkeep_T_108,_xbar_level0_io_s_axis_tkeep_T_107,
    _xbar_level0_io_s_axis_tkeep_T_106,_xbar_level0_io_s_axis_tkeep_T_105,_xbar_level0_io_s_axis_tkeep_T_104,
    xbar_level0_io_s_axis_tkeep_hi_lo_lo}; // @[bfs_remote.scala 654:124]
  wire [7:0] xbar_level0_io_s_axis_tkeep_hi_hi_lo = {_xbar_level0_io_s_axis_tkeep_T_119,
    _xbar_level0_io_s_axis_tkeep_T_118,_xbar_level0_io_s_axis_tkeep_T_117,_xbar_level0_io_s_axis_tkeep_T_116,
    _xbar_level0_io_s_axis_tkeep_T_115,_xbar_level0_io_s_axis_tkeep_T_114,_xbar_level0_io_s_axis_tkeep_T_113,
    _xbar_level0_io_s_axis_tkeep_T_112}; // @[bfs_remote.scala 654:124]
  wire [31:0] xbar_level0_io_s_axis_tkeep_hi = {_xbar_level0_io_s_axis_tkeep_T_127,_xbar_level0_io_s_axis_tkeep_T_126,
    _xbar_level0_io_s_axis_tkeep_T_125,_xbar_level0_io_s_axis_tkeep_T_124,_xbar_level0_io_s_axis_tkeep_T_123,
    _xbar_level0_io_s_axis_tkeep_T_122,_xbar_level0_io_s_axis_tkeep_T_121,_xbar_level0_io_s_axis_tkeep_T_120,
    xbar_level0_io_s_axis_tkeep_hi_hi_lo,xbar_level0_io_s_axis_tkeep_hi_lo}; // @[bfs_remote.scala 654:124]
  wire  _filtered_keep_0_T_4 = xbar_level0_m_axis_tdata[1:0] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_0_T_5 = xbar_level0_m_axis_tdata[31] | _filtered_keep_0_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_0 = xbar_level0_m_axis_tkeep[0] & _filtered_keep_0_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_1_T_4 = xbar_level0_m_axis_tdata[33:32] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_1_T_5 = xbar_level0_m_axis_tdata[63] | _filtered_keep_1_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_1 = xbar_level0_m_axis_tkeep[1] & _filtered_keep_1_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_2_T_4 = xbar_level0_m_axis_tdata[65:64] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_2_T_5 = xbar_level0_m_axis_tdata[95] | _filtered_keep_2_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_2 = xbar_level0_m_axis_tkeep[2] & _filtered_keep_2_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_3_T_4 = xbar_level0_m_axis_tdata[97:96] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_3_T_5 = xbar_level0_m_axis_tdata[127] | _filtered_keep_3_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_3 = xbar_level0_m_axis_tkeep[3] & _filtered_keep_3_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_4_T_4 = xbar_level0_m_axis_tdata[129:128] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_4_T_5 = xbar_level0_m_axis_tdata[159] | _filtered_keep_4_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_4 = xbar_level0_m_axis_tkeep[4] & _filtered_keep_4_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_5_T_4 = xbar_level0_m_axis_tdata[161:160] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_5_T_5 = xbar_level0_m_axis_tdata[191] | _filtered_keep_5_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_5 = xbar_level0_m_axis_tkeep[5] & _filtered_keep_5_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_6_T_4 = xbar_level0_m_axis_tdata[193:192] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_6_T_5 = xbar_level0_m_axis_tdata[223] | _filtered_keep_6_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_6 = xbar_level0_m_axis_tkeep[6] & _filtered_keep_6_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_7_T_4 = xbar_level0_m_axis_tdata[225:224] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_7_T_5 = xbar_level0_m_axis_tdata[255] | _filtered_keep_7_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_7 = xbar_level0_m_axis_tkeep[7] & _filtered_keep_7_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_8_T_4 = xbar_level0_m_axis_tdata[257:256] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_8_T_5 = xbar_level0_m_axis_tdata[287] | _filtered_keep_8_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_8 = xbar_level0_m_axis_tkeep[8] & _filtered_keep_8_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_9_T_4 = xbar_level0_m_axis_tdata[289:288] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_9_T_5 = xbar_level0_m_axis_tdata[319] | _filtered_keep_9_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_9 = xbar_level0_m_axis_tkeep[9] & _filtered_keep_9_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_10_T_4 = xbar_level0_m_axis_tdata[321:320] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_10_T_5 = xbar_level0_m_axis_tdata[351] | _filtered_keep_10_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_10 = xbar_level0_m_axis_tkeep[10] & _filtered_keep_10_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_11_T_4 = xbar_level0_m_axis_tdata[353:352] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_11_T_5 = xbar_level0_m_axis_tdata[383] | _filtered_keep_11_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_11 = xbar_level0_m_axis_tkeep[11] & _filtered_keep_11_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_12_T_4 = xbar_level0_m_axis_tdata[385:384] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_12_T_5 = xbar_level0_m_axis_tdata[415] | _filtered_keep_12_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_12 = xbar_level0_m_axis_tkeep[12] & _filtered_keep_12_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_13_T_4 = xbar_level0_m_axis_tdata[417:416] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_13_T_5 = xbar_level0_m_axis_tdata[447] | _filtered_keep_13_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_13 = xbar_level0_m_axis_tkeep[13] & _filtered_keep_13_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_14_T_4 = xbar_level0_m_axis_tdata[449:448] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_14_T_5 = xbar_level0_m_axis_tdata[479] | _filtered_keep_14_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_14 = xbar_level0_m_axis_tkeep[14] & _filtered_keep_14_T_5; // @[bfs_remote.scala 670:15]
  wire  _filtered_keep_15_T_4 = xbar_level0_m_axis_tdata[481:480] == local_fpga_id; // @[bfs_remote.scala 664:36]
  wire  _filtered_keep_15_T_5 = xbar_level0_m_axis_tdata[511] | _filtered_keep_15_T_4; // @[bfs_remote.scala 671:12]
  wire  filtered_keep_15 = xbar_level0_m_axis_tkeep[15] & _filtered_keep_15_T_5; // @[bfs_remote.scala 670:15]
  reg  flush_reg; // @[bfs_remote.scala 676:26]
  wire  _GEN_0 = io_flush | flush_reg; // @[bfs_remote.scala 679:23 bfs_remote.scala 680:15 bfs_remote.scala 676:26]
  wire [7:0] collector_io_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[bfs_remote.scala 684:53]
  wire [7:0] collector_io_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[bfs_remote.scala 684:53]
  wire [3:0] xbar_level0_io_m_axis_tready_hi_1 = {io_remote_out_3_ready,io_remote_out_2_ready,io_remote_out_1_ready,
    io_remote_out_0_ready}; // @[bfs_remote.scala 687:84]
  wire [511:0] _in_data_WIRE = switch_level1_io_out_bits_tdata;
  wire [31:0] in_data_0 = _in_data_WIRE[31:0]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_1 = _in_data_WIRE[63:32]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_2 = _in_data_WIRE[95:64]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_3 = _in_data_WIRE[127:96]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_4 = _in_data_WIRE[159:128]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_5 = _in_data_WIRE[191:160]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_6 = _in_data_WIRE[223:192]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_7 = _in_data_WIRE[255:224]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_8 = _in_data_WIRE[287:256]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_9 = _in_data_WIRE[319:288]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_10 = _in_data_WIRE[351:320]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_11 = _in_data_WIRE[383:352]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_12 = _in_data_WIRE[415:384]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_13 = _in_data_WIRE[447:416]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_14 = _in_data_WIRE[479:448]; // @[bfs_remote.scala 713:57]
  wire [31:0] in_data_15 = _in_data_WIRE[511:480]; // @[bfs_remote.scala 713:57]
  wire  in_keep_0 = switch_level1_io_out_bits_tkeep[0]; // @[bfs_remote.scala 714:71]
  wire  in_keep_1 = switch_level1_io_out_bits_tkeep[1]; // @[bfs_remote.scala 714:71]
  wire  in_keep_2 = switch_level1_io_out_bits_tkeep[2]; // @[bfs_remote.scala 714:71]
  wire  in_keep_3 = switch_level1_io_out_bits_tkeep[3]; // @[bfs_remote.scala 714:71]
  wire  in_keep_4 = switch_level1_io_out_bits_tkeep[4]; // @[bfs_remote.scala 714:71]
  wire  in_keep_5 = switch_level1_io_out_bits_tkeep[5]; // @[bfs_remote.scala 714:71]
  wire  in_keep_6 = switch_level1_io_out_bits_tkeep[6]; // @[bfs_remote.scala 714:71]
  wire  in_keep_7 = switch_level1_io_out_bits_tkeep[7]; // @[bfs_remote.scala 714:71]
  wire  in_keep_8 = switch_level1_io_out_bits_tkeep[8]; // @[bfs_remote.scala 714:71]
  wire  in_keep_9 = switch_level1_io_out_bits_tkeep[9]; // @[bfs_remote.scala 714:71]
  wire  in_keep_10 = switch_level1_io_out_bits_tkeep[10]; // @[bfs_remote.scala 714:71]
  wire  in_keep_11 = switch_level1_io_out_bits_tkeep[11]; // @[bfs_remote.scala 714:71]
  wire  in_keep_12 = switch_level1_io_out_bits_tkeep[12]; // @[bfs_remote.scala 714:71]
  wire  in_keep_13 = switch_level1_io_out_bits_tkeep[13]; // @[bfs_remote.scala 714:71]
  wire  in_keep_14 = switch_level1_io_out_bits_tkeep[14]; // @[bfs_remote.scala 714:71]
  wire  replication_1 = in_data_0 == in_data_1 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_2_T_1 = in_data_0 == in_data_2 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_2_T_3 = in_data_1 == in_data_2 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  replication_2 = _replication_2_T_1 | _replication_2_T_3; // @[bfs_remote.scala 721:17]
  wire  _replication_3_T_1 = in_data_0 == in_data_3 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_3_T_3 = in_data_1 == in_data_3 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_3_T_5 = in_data_2 == in_data_3 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  replication_3 = _replication_3_T_1 | _replication_3_T_3 | _replication_3_T_5; // @[bfs_remote.scala 721:17]
  wire  _replication_4_T_1 = in_data_0 == in_data_4 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_4_T_3 = in_data_1 == in_data_4 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_4_T_5 = in_data_2 == in_data_4 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_4_T_7 = in_data_3 == in_data_4 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  replication_4 = _replication_4_T_1 | _replication_4_T_3 | _replication_4_T_5 | _replication_4_T_7; // @[bfs_remote.scala 721:17]
  wire  _replication_5_T_1 = in_data_0 == in_data_5 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_5_T_3 = in_data_1 == in_data_5 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_5_T_5 = in_data_2 == in_data_5 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_5_T_7 = in_data_3 == in_data_5 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_5_T_9 = in_data_4 == in_data_5 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  replication_5 = _replication_5_T_1 | _replication_5_T_3 | _replication_5_T_5 | _replication_5_T_7 |
    _replication_5_T_9; // @[bfs_remote.scala 721:17]
  wire  _replication_6_T_1 = in_data_0 == in_data_6 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_6_T_3 = in_data_1 == in_data_6 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_6_T_5 = in_data_2 == in_data_6 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_6_T_7 = in_data_3 == in_data_6 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_6_T_9 = in_data_4 == in_data_6 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_6_T_11 = in_data_5 == in_data_6 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  replication_6 = _replication_6_T_1 | _replication_6_T_3 | _replication_6_T_5 | _replication_6_T_7 |
    _replication_6_T_9 | _replication_6_T_11; // @[bfs_remote.scala 721:17]
  wire  _replication_7_T_1 = in_data_0 == in_data_7 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_7_T_3 = in_data_1 == in_data_7 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_7_T_5 = in_data_2 == in_data_7 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_7_T_7 = in_data_3 == in_data_7 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_7_T_9 = in_data_4 == in_data_7 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_7_T_11 = in_data_5 == in_data_7 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  _replication_7_T_13 = in_data_6 == in_data_7 & in_keep_6; // @[bfs_remote.scala 720:47]
  wire  replication_7 = _replication_7_T_1 | _replication_7_T_3 | _replication_7_T_5 | _replication_7_T_7 |
    _replication_7_T_9 | _replication_7_T_11 | _replication_7_T_13; // @[bfs_remote.scala 721:17]
  wire  _replication_8_T_1 = in_data_0 == in_data_8 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_8_T_3 = in_data_1 == in_data_8 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_8_T_5 = in_data_2 == in_data_8 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_8_T_7 = in_data_3 == in_data_8 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_8_T_9 = in_data_4 == in_data_8 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_8_T_11 = in_data_5 == in_data_8 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  _replication_8_T_13 = in_data_6 == in_data_8 & in_keep_6; // @[bfs_remote.scala 720:47]
  wire  _replication_8_T_15 = in_data_7 == in_data_8 & in_keep_7; // @[bfs_remote.scala 720:47]
  wire  replication_8 = _replication_8_T_1 | _replication_8_T_3 | _replication_8_T_5 | _replication_8_T_7 |
    _replication_8_T_9 | _replication_8_T_11 | _replication_8_T_13 | _replication_8_T_15; // @[bfs_remote.scala 721:17]
  wire  _replication_9_T_1 = in_data_0 == in_data_9 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_9_T_3 = in_data_1 == in_data_9 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_9_T_5 = in_data_2 == in_data_9 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_9_T_7 = in_data_3 == in_data_9 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_9_T_9 = in_data_4 == in_data_9 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_9_T_11 = in_data_5 == in_data_9 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  _replication_9_T_13 = in_data_6 == in_data_9 & in_keep_6; // @[bfs_remote.scala 720:47]
  wire  _replication_9_T_15 = in_data_7 == in_data_9 & in_keep_7; // @[bfs_remote.scala 720:47]
  wire  _replication_9_T_17 = in_data_8 == in_data_9 & in_keep_8; // @[bfs_remote.scala 720:47]
  wire  replication_9 = _replication_9_T_1 | _replication_9_T_3 | _replication_9_T_5 | _replication_9_T_7 |
    _replication_9_T_9 | _replication_9_T_11 | _replication_9_T_13 | _replication_9_T_15 | _replication_9_T_17; // @[bfs_remote.scala 721:17]
  wire  _replication_10_T_1 = in_data_0 == in_data_10 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_10_T_3 = in_data_1 == in_data_10 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_10_T_5 = in_data_2 == in_data_10 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_10_T_7 = in_data_3 == in_data_10 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_10_T_9 = in_data_4 == in_data_10 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_10_T_11 = in_data_5 == in_data_10 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  _replication_10_T_13 = in_data_6 == in_data_10 & in_keep_6; // @[bfs_remote.scala 720:47]
  wire  _replication_10_T_15 = in_data_7 == in_data_10 & in_keep_7; // @[bfs_remote.scala 720:47]
  wire  _replication_10_T_17 = in_data_8 == in_data_10 & in_keep_8; // @[bfs_remote.scala 720:47]
  wire  _replication_10_T_19 = in_data_9 == in_data_10 & in_keep_9; // @[bfs_remote.scala 720:47]
  wire  replication_10 = _replication_10_T_1 | _replication_10_T_3 | _replication_10_T_5 | _replication_10_T_7 |
    _replication_10_T_9 | _replication_10_T_11 | _replication_10_T_13 | _replication_10_T_15 | _replication_10_T_17 |
    _replication_10_T_19; // @[bfs_remote.scala 721:17]
  wire  _replication_11_T_1 = in_data_0 == in_data_11 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_3 = in_data_1 == in_data_11 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_5 = in_data_2 == in_data_11 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_7 = in_data_3 == in_data_11 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_9 = in_data_4 == in_data_11 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_11 = in_data_5 == in_data_11 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_13 = in_data_6 == in_data_11 & in_keep_6; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_15 = in_data_7 == in_data_11 & in_keep_7; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_17 = in_data_8 == in_data_11 & in_keep_8; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_19 = in_data_9 == in_data_11 & in_keep_9; // @[bfs_remote.scala 720:47]
  wire  _replication_11_T_21 = in_data_10 == in_data_11 & in_keep_10; // @[bfs_remote.scala 720:47]
  wire  replication_11 = _replication_11_T_1 | _replication_11_T_3 | _replication_11_T_5 | _replication_11_T_7 |
    _replication_11_T_9 | _replication_11_T_11 | _replication_11_T_13 | _replication_11_T_15 | _replication_11_T_17 |
    _replication_11_T_19 | _replication_11_T_21; // @[bfs_remote.scala 721:17]
  wire  _replication_12_T_1 = in_data_0 == in_data_12 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_3 = in_data_1 == in_data_12 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_5 = in_data_2 == in_data_12 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_7 = in_data_3 == in_data_12 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_9 = in_data_4 == in_data_12 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_11 = in_data_5 == in_data_12 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_13 = in_data_6 == in_data_12 & in_keep_6; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_15 = in_data_7 == in_data_12 & in_keep_7; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_17 = in_data_8 == in_data_12 & in_keep_8; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_19 = in_data_9 == in_data_12 & in_keep_9; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_21 = in_data_10 == in_data_12 & in_keep_10; // @[bfs_remote.scala 720:47]
  wire  _replication_12_T_23 = in_data_11 == in_data_12 & in_keep_11; // @[bfs_remote.scala 720:47]
  wire  replication_12 = _replication_12_T_1 | _replication_12_T_3 | _replication_12_T_5 | _replication_12_T_7 |
    _replication_12_T_9 | _replication_12_T_11 | _replication_12_T_13 | _replication_12_T_15 | _replication_12_T_17 |
    _replication_12_T_19 | _replication_12_T_21 | _replication_12_T_23; // @[bfs_remote.scala 721:17]
  wire  _replication_13_T_1 = in_data_0 == in_data_13 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_3 = in_data_1 == in_data_13 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_5 = in_data_2 == in_data_13 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_7 = in_data_3 == in_data_13 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_9 = in_data_4 == in_data_13 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_11 = in_data_5 == in_data_13 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_13 = in_data_6 == in_data_13 & in_keep_6; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_15 = in_data_7 == in_data_13 & in_keep_7; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_17 = in_data_8 == in_data_13 & in_keep_8; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_19 = in_data_9 == in_data_13 & in_keep_9; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_21 = in_data_10 == in_data_13 & in_keep_10; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_23 = in_data_11 == in_data_13 & in_keep_11; // @[bfs_remote.scala 720:47]
  wire  _replication_13_T_25 = in_data_12 == in_data_13 & in_keep_12; // @[bfs_remote.scala 720:47]
  wire  replication_13 = _replication_13_T_1 | _replication_13_T_3 | _replication_13_T_5 | _replication_13_T_7 |
    _replication_13_T_9 | _replication_13_T_11 | _replication_13_T_13 | _replication_13_T_15 | _replication_13_T_17 |
    _replication_13_T_19 | _replication_13_T_21 | _replication_13_T_23 | _replication_13_T_25; // @[bfs_remote.scala 721:17]
  wire  _replication_14_T_1 = in_data_0 == in_data_14 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_3 = in_data_1 == in_data_14 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_5 = in_data_2 == in_data_14 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_7 = in_data_3 == in_data_14 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_9 = in_data_4 == in_data_14 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_11 = in_data_5 == in_data_14 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_13 = in_data_6 == in_data_14 & in_keep_6; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_15 = in_data_7 == in_data_14 & in_keep_7; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_17 = in_data_8 == in_data_14 & in_keep_8; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_19 = in_data_9 == in_data_14 & in_keep_9; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_21 = in_data_10 == in_data_14 & in_keep_10; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_23 = in_data_11 == in_data_14 & in_keep_11; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_25 = in_data_12 == in_data_14 & in_keep_12; // @[bfs_remote.scala 720:47]
  wire  _replication_14_T_27 = in_data_13 == in_data_14 & in_keep_13; // @[bfs_remote.scala 720:47]
  wire  replication_14 = _replication_14_T_1 | _replication_14_T_3 | _replication_14_T_5 | _replication_14_T_7 |
    _replication_14_T_9 | _replication_14_T_11 | _replication_14_T_13 | _replication_14_T_15 | _replication_14_T_17 |
    _replication_14_T_19 | _replication_14_T_21 | _replication_14_T_23 | _replication_14_T_25 | _replication_14_T_27; // @[bfs_remote.scala 721:17]
  wire  _replication_15_T_1 = in_data_0 == in_data_15 & in_keep_0; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_3 = in_data_1 == in_data_15 & in_keep_1; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_5 = in_data_2 == in_data_15 & in_keep_2; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_7 = in_data_3 == in_data_15 & in_keep_3; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_9 = in_data_4 == in_data_15 & in_keep_4; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_11 = in_data_5 == in_data_15 & in_keep_5; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_13 = in_data_6 == in_data_15 & in_keep_6; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_15 = in_data_7 == in_data_15 & in_keep_7; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_17 = in_data_8 == in_data_15 & in_keep_8; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_19 = in_data_9 == in_data_15 & in_keep_9; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_21 = in_data_10 == in_data_15 & in_keep_10; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_23 = in_data_11 == in_data_15 & in_keep_11; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_25 = in_data_12 == in_data_15 & in_keep_12; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_27 = in_data_13 == in_data_15 & in_keep_13; // @[bfs_remote.scala 720:47]
  wire  _replication_15_T_29 = in_data_14 == in_data_15 & in_keep_14; // @[bfs_remote.scala 720:47]
  wire  replication_15 = _replication_15_T_1 | _replication_15_T_3 | _replication_15_T_5 | _replication_15_T_7 |
    _replication_15_T_9 | _replication_15_T_11 | _replication_15_T_13 | _replication_15_T_15 | _replication_15_T_17 |
    _replication_15_T_19 | _replication_15_T_21 | _replication_15_T_23 | _replication_15_T_25 | _replication_15_T_27 |
    _replication_15_T_29; // @[bfs_remote.scala 721:17]
  wire  _mid_io_s_axis_tkeep_T_1 = ~replication_1; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_2 = ~replication_2; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_3 = ~replication_3; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_4 = ~replication_4; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_5 = ~replication_5; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_6 = ~replication_6; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_7 = ~replication_7; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_8 = ~replication_8; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_9 = ~replication_9; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_10 = ~replication_10; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_11 = ~replication_11; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_12 = ~replication_12; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_13 = ~replication_13; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_14 = ~replication_14; // @[bfs_remote.scala 730:84]
  wire  _mid_io_s_axis_tkeep_T_15 = ~replication_15; // @[bfs_remote.scala 730:84]
  wire [7:0] mid_io_s_axis_tkeep_lo = {_mid_io_s_axis_tkeep_T_7,_mid_io_s_axis_tkeep_T_6,_mid_io_s_axis_tkeep_T_5,
    _mid_io_s_axis_tkeep_T_4,_mid_io_s_axis_tkeep_T_3,_mid_io_s_axis_tkeep_T_2,_mid_io_s_axis_tkeep_T_1,1'h1}; // @[bfs_remote.scala 730:95]
  wire [15:0] _mid_io_s_axis_tkeep_T_16 = {_mid_io_s_axis_tkeep_T_15,_mid_io_s_axis_tkeep_T_14,_mid_io_s_axis_tkeep_T_13
    ,_mid_io_s_axis_tkeep_T_12,_mid_io_s_axis_tkeep_T_11,_mid_io_s_axis_tkeep_T_10,_mid_io_s_axis_tkeep_T_9,
    _mid_io_s_axis_tkeep_T_8,mid_io_s_axis_tkeep_lo}; // @[bfs_remote.scala 730:95]
  wire [63:0] _GEN_2 = {{48'd0}, _mid_io_s_axis_tkeep_T_16}; // @[bfs_remote.scala 730:58]
  wire  _xbar_level1_io_s_axis_tkeep_T_64 = mid_m_axis_tkeep[0] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_65 = mid_m_axis_tkeep[1] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_66 = mid_m_axis_tkeep[2] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_67 = mid_m_axis_tkeep[3] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_68 = mid_m_axis_tkeep[4] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_69 = mid_m_axis_tkeep[5] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_70 = mid_m_axis_tkeep[6] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_71 = mid_m_axis_tkeep[7] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_72 = mid_m_axis_tkeep[8] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_73 = mid_m_axis_tkeep[9] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_74 = mid_m_axis_tkeep[10] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_75 = mid_m_axis_tkeep[11] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_76 = mid_m_axis_tkeep[12] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_77 = mid_m_axis_tkeep[13] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_78 = mid_m_axis_tkeep[14] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_79 = mid_m_axis_tkeep[15] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_80 = mid_m_axis_tkeep[16] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_81 = mid_m_axis_tkeep[17] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_82 = mid_m_axis_tkeep[18] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_83 = mid_m_axis_tkeep[19] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_84 = mid_m_axis_tkeep[20] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_85 = mid_m_axis_tkeep[21] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_86 = mid_m_axis_tkeep[22] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_87 = mid_m_axis_tkeep[23] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_88 = mid_m_axis_tkeep[24] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_89 = mid_m_axis_tkeep[25] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_90 = mid_m_axis_tkeep[26] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_91 = mid_m_axis_tkeep[27] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_92 = mid_m_axis_tkeep[28] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_93 = mid_m_axis_tkeep[29] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_94 = mid_m_axis_tkeep[30] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_95 = mid_m_axis_tkeep[31] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_96 = mid_m_axis_tkeep[32] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_97 = mid_m_axis_tkeep[33] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_98 = mid_m_axis_tkeep[34] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_99 = mid_m_axis_tkeep[35] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_100 = mid_m_axis_tkeep[36] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_101 = mid_m_axis_tkeep[37] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_102 = mid_m_axis_tkeep[38] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_103 = mid_m_axis_tkeep[39] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_104 = mid_m_axis_tkeep[40] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_105 = mid_m_axis_tkeep[41] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_106 = mid_m_axis_tkeep[42] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_107 = mid_m_axis_tkeep[43] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_108 = mid_m_axis_tkeep[44] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_109 = mid_m_axis_tkeep[45] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_110 = mid_m_axis_tkeep[46] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_111 = mid_m_axis_tkeep[47] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_112 = mid_m_axis_tkeep[48] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_113 = mid_m_axis_tkeep[49] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_114 = mid_m_axis_tkeep[50] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_115 = mid_m_axis_tkeep[51] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_116 = mid_m_axis_tkeep[52] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_117 = mid_m_axis_tkeep[53] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_118 = mid_m_axis_tkeep[54] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_119 = mid_m_axis_tkeep[55] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_120 = mid_m_axis_tkeep[56] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_121 = mid_m_axis_tkeep[57] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_122 = mid_m_axis_tkeep[58] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_123 = mid_m_axis_tkeep[59] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_124 = mid_m_axis_tkeep[60] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_125 = mid_m_axis_tkeep[61] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_126 = mid_m_axis_tkeep[62] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire  _xbar_level1_io_s_axis_tkeep_T_127 = mid_m_axis_tkeep[63] & mid_m_axis_tvalid; // @[bfs_remote.scala 738:83]
  wire [7:0] xbar_level1_io_s_axis_tkeep_lo_lo_lo = {_xbar_level1_io_s_axis_tkeep_T_71,_xbar_level1_io_s_axis_tkeep_T_70
    ,_xbar_level1_io_s_axis_tkeep_T_69,_xbar_level1_io_s_axis_tkeep_T_68,_xbar_level1_io_s_axis_tkeep_T_67,
    _xbar_level1_io_s_axis_tkeep_T_66,_xbar_level1_io_s_axis_tkeep_T_65,_xbar_level1_io_s_axis_tkeep_T_64}; // @[bfs_remote.scala 738:114]
  wire [15:0] xbar_level1_io_s_axis_tkeep_lo_lo = {_xbar_level1_io_s_axis_tkeep_T_79,_xbar_level1_io_s_axis_tkeep_T_78,
    _xbar_level1_io_s_axis_tkeep_T_77,_xbar_level1_io_s_axis_tkeep_T_76,_xbar_level1_io_s_axis_tkeep_T_75,
    _xbar_level1_io_s_axis_tkeep_T_74,_xbar_level1_io_s_axis_tkeep_T_73,_xbar_level1_io_s_axis_tkeep_T_72,
    xbar_level1_io_s_axis_tkeep_lo_lo_lo}; // @[bfs_remote.scala 738:114]
  wire [7:0] xbar_level1_io_s_axis_tkeep_lo_hi_lo = {_xbar_level1_io_s_axis_tkeep_T_87,_xbar_level1_io_s_axis_tkeep_T_86
    ,_xbar_level1_io_s_axis_tkeep_T_85,_xbar_level1_io_s_axis_tkeep_T_84,_xbar_level1_io_s_axis_tkeep_T_83,
    _xbar_level1_io_s_axis_tkeep_T_82,_xbar_level1_io_s_axis_tkeep_T_81,_xbar_level1_io_s_axis_tkeep_T_80}; // @[bfs_remote.scala 738:114]
  wire [31:0] xbar_level1_io_s_axis_tkeep_lo = {_xbar_level1_io_s_axis_tkeep_T_95,_xbar_level1_io_s_axis_tkeep_T_94,
    _xbar_level1_io_s_axis_tkeep_T_93,_xbar_level1_io_s_axis_tkeep_T_92,_xbar_level1_io_s_axis_tkeep_T_91,
    _xbar_level1_io_s_axis_tkeep_T_90,_xbar_level1_io_s_axis_tkeep_T_89,_xbar_level1_io_s_axis_tkeep_T_88,
    xbar_level1_io_s_axis_tkeep_lo_hi_lo,xbar_level1_io_s_axis_tkeep_lo_lo}; // @[bfs_remote.scala 738:114]
  wire [7:0] xbar_level1_io_s_axis_tkeep_hi_lo_lo = {_xbar_level1_io_s_axis_tkeep_T_103,
    _xbar_level1_io_s_axis_tkeep_T_102,_xbar_level1_io_s_axis_tkeep_T_101,_xbar_level1_io_s_axis_tkeep_T_100,
    _xbar_level1_io_s_axis_tkeep_T_99,_xbar_level1_io_s_axis_tkeep_T_98,_xbar_level1_io_s_axis_tkeep_T_97,
    _xbar_level1_io_s_axis_tkeep_T_96}; // @[bfs_remote.scala 738:114]
  wire [15:0] xbar_level1_io_s_axis_tkeep_hi_lo = {_xbar_level1_io_s_axis_tkeep_T_111,_xbar_level1_io_s_axis_tkeep_T_110
    ,_xbar_level1_io_s_axis_tkeep_T_109,_xbar_level1_io_s_axis_tkeep_T_108,_xbar_level1_io_s_axis_tkeep_T_107,
    _xbar_level1_io_s_axis_tkeep_T_106,_xbar_level1_io_s_axis_tkeep_T_105,_xbar_level1_io_s_axis_tkeep_T_104,
    xbar_level1_io_s_axis_tkeep_hi_lo_lo}; // @[bfs_remote.scala 738:114]
  wire [7:0] xbar_level1_io_s_axis_tkeep_hi_hi_lo = {_xbar_level1_io_s_axis_tkeep_T_119,
    _xbar_level1_io_s_axis_tkeep_T_118,_xbar_level1_io_s_axis_tkeep_T_117,_xbar_level1_io_s_axis_tkeep_T_116,
    _xbar_level1_io_s_axis_tkeep_T_115,_xbar_level1_io_s_axis_tkeep_T_114,_xbar_level1_io_s_axis_tkeep_T_113,
    _xbar_level1_io_s_axis_tkeep_T_112}; // @[bfs_remote.scala 738:114]
  wire [31:0] xbar_level1_io_s_axis_tkeep_hi = {_xbar_level1_io_s_axis_tkeep_T_127,_xbar_level1_io_s_axis_tkeep_T_126,
    _xbar_level1_io_s_axis_tkeep_T_125,_xbar_level1_io_s_axis_tkeep_T_124,_xbar_level1_io_s_axis_tkeep_T_123,
    _xbar_level1_io_s_axis_tkeep_T_122,_xbar_level1_io_s_axis_tkeep_T_121,_xbar_level1_io_s_axis_tkeep_T_120,
    xbar_level1_io_s_axis_tkeep_hi_hi_lo,xbar_level1_io_s_axis_tkeep_hi_lo}; // @[bfs_remote.scala 738:114]
  wire  _xbar_level1_io_m_axis_tready_WIRE_1 = backend_1_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_0 = backend_0_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_3 = backend_3_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_2 = backend_2_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_5 = backend_5_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_4 = backend_4_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_7 = backend_7_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_6 = backend_6_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire [7:0] xbar_level1_io_m_axis_tready_lo = {_xbar_level1_io_m_axis_tready_WIRE_7,
    _xbar_level1_io_m_axis_tready_WIRE_6,_xbar_level1_io_m_axis_tready_WIRE_5,_xbar_level1_io_m_axis_tready_WIRE_4,
    _xbar_level1_io_m_axis_tready_WIRE_3,_xbar_level1_io_m_axis_tready_WIRE_2,_xbar_level1_io_m_axis_tready_WIRE_1,
    _xbar_level1_io_m_axis_tready_WIRE_0}; // @[bfs_remote.scala 754:12]
  wire  _xbar_level1_io_m_axis_tready_WIRE_9 = backend_9_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_8 = backend_8_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_11 = backend_11_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_10 = backend_10_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_13 = backend_13_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_12 = backend_12_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_15 = backend_15_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire  _xbar_level1_io_m_axis_tready_WIRE_14 = backend_14_s_axis_tready; // @[bfs_remote.scala 752:63 bfs_remote.scala 752:63]
  wire [7:0] xbar_level1_io_m_axis_tready_hi = {_xbar_level1_io_m_axis_tready_WIRE_15,
    _xbar_level1_io_m_axis_tready_WIRE_14,_xbar_level1_io_m_axis_tready_WIRE_13,_xbar_level1_io_m_axis_tready_WIRE_12,
    _xbar_level1_io_m_axis_tready_WIRE_11,_xbar_level1_io_m_axis_tready_WIRE_10,_xbar_level1_io_m_axis_tready_WIRE_9,
    _xbar_level1_io_m_axis_tready_WIRE_8}; // @[bfs_remote.scala 754:12]
  wire [63:0] _io_pe_out_0_bits_tkeep_T = backend_0_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_1_bits_tkeep_T = backend_1_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_2_bits_tkeep_T = backend_2_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_3_bits_tkeep_T = backend_3_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_4_bits_tkeep_T = backend_4_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_5_bits_tkeep_T = backend_5_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_6_bits_tkeep_T = backend_6_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_7_bits_tkeep_T = backend_7_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_8_bits_tkeep_T = backend_8_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_9_bits_tkeep_T = backend_9_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_10_bits_tkeep_T = backend_10_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_11_bits_tkeep_T = backend_11_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_12_bits_tkeep_T = backend_12_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_13_bits_tkeep_T = backend_13_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_14_bits_tkeep_T = backend_14_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  wire [63:0] _io_pe_out_15_bits_tkeep_T = backend_15_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  axis_combiner_level0 combiner_level0 ( // @[bfs_remote.scala 628:31]
    .aclk(combiner_level0_aclk),
    .aresetn(combiner_level0_aresetn),
    .s_axis_tdata(combiner_level0_s_axis_tdata),
    .s_axis_tvalid(combiner_level0_s_axis_tvalid),
    .s_axis_tkeep(combiner_level0_s_axis_tkeep),
    .s_axis_tready(combiner_level0_s_axis_tready),
    .s_axis_tlast(combiner_level0_s_axis_tlast),
    .s_axis_tid(combiner_level0_s_axis_tid),
    .m_axis_tdata(combiner_level0_m_axis_tdata),
    .m_axis_tvalid(combiner_level0_m_axis_tvalid),
    .m_axis_tkeep(combiner_level0_m_axis_tkeep),
    .m_axis_tready(combiner_level0_m_axis_tready),
    .m_axis_tlast(combiner_level0_m_axis_tlast),
    .m_axis_tid(combiner_level0_m_axis_tid)
  );
  Remote_xbar_reg_slice frontend ( // @[bfs_remote.scala 640:24]
    .aclk(frontend_aclk),
    .aresetn(frontend_aresetn),
    .s_axis_tdata(frontend_s_axis_tdata),
    .s_axis_tvalid(frontend_s_axis_tvalid),
    .s_axis_tkeep(frontend_s_axis_tkeep),
    .s_axis_tready(frontend_s_axis_tready),
    .s_axis_tlast(frontend_s_axis_tlast),
    .m_axis_tdata(frontend_m_axis_tdata),
    .m_axis_tvalid(frontend_m_axis_tvalid),
    .m_axis_tkeep(frontend_m_axis_tkeep),
    .m_axis_tready(frontend_m_axis_tready),
    .m_axis_tlast(frontend_m_axis_tlast)
  );
  axis_broadcaster_level0 xbar_level0 ( // @[bfs_remote.scala 649:27]
    .aclk(xbar_level0_aclk),
    .aresetn(xbar_level0_aresetn),
    .s_axis_tdata(xbar_level0_s_axis_tdata),
    .s_axis_tvalid(xbar_level0_s_axis_tvalid),
    .s_axis_tkeep(xbar_level0_s_axis_tkeep),
    .s_axis_tready(xbar_level0_s_axis_tready),
    .s_axis_tlast(xbar_level0_s_axis_tlast),
    .s_axis_tid(xbar_level0_s_axis_tid),
    .m_axis_tdata(xbar_level0_m_axis_tdata),
    .m_axis_tvalid(xbar_level0_m_axis_tvalid),
    .m_axis_tkeep(xbar_level0_m_axis_tkeep),
    .m_axis_tready(xbar_level0_m_axis_tready),
    .m_axis_tlast(xbar_level0_m_axis_tlast),
    .m_axis_tid(xbar_level0_m_axis_tid)
  );
  axis_data_collector collector ( // @[bfs_remote.scala 682:25]
    .clock(collector_clock),
    .reset(collector_reset),
    .io_in_ready(collector_io_in_ready),
    .io_in_valid(collector_io_in_valid),
    .io_in_bits_tdata(collector_io_in_bits_tdata),
    .io_in_bits_tkeep(collector_io_in_bits_tkeep),
    .io_out_ready(collector_io_out_ready),
    .io_out_valid(collector_io_out_valid),
    .io_out_bits_tdata(collector_io_out_bits_tdata),
    .io_out_bits_tkeep(collector_io_out_bits_tkeep),
    .io_out_bits_tlast(collector_io_out_bits_tlast),
    .io_flush(collector_io_flush),
    .io_empty(collector_io_empty)
  );
  Remote_xbar_buffer1 buffer1 ( // @[bfs_remote.scala 690:23]
    .s_axis_aclk(buffer1_s_axis_aclk),
    .s_axis_aresetn(buffer1_s_axis_aresetn),
    .s_axis_tdata(buffer1_s_axis_tdata),
    .s_axis_tvalid(buffer1_s_axis_tvalid),
    .s_axis_tkeep(buffer1_s_axis_tkeep),
    .s_axis_tready(buffer1_s_axis_tready),
    .s_axis_tlast(buffer1_s_axis_tlast),
    .s_axis_tid(buffer1_s_axis_tid),
    .m_axis_tdata(buffer1_m_axis_tdata),
    .m_axis_tvalid(buffer1_m_axis_tvalid),
    .m_axis_tkeep(buffer1_m_axis_tkeep),
    .m_axis_tready(buffer1_m_axis_tready),
    .m_axis_tlast(buffer1_m_axis_tlast),
    .m_axis_tid(buffer1_m_axis_tid)
  );
  Remote_xbar_reg_slice remote_in_reg ( // @[bfs_remote.scala 697:29]
    .aclk(remote_in_reg_aclk),
    .aresetn(remote_in_reg_aresetn),
    .s_axis_tdata(remote_in_reg_s_axis_tdata),
    .s_axis_tvalid(remote_in_reg_s_axis_tvalid),
    .s_axis_tkeep(remote_in_reg_s_axis_tkeep),
    .s_axis_tready(remote_in_reg_s_axis_tready),
    .s_axis_tlast(remote_in_reg_s_axis_tlast),
    .m_axis_tdata(remote_in_reg_m_axis_tdata),
    .m_axis_tvalid(remote_in_reg_m_axis_tvalid),
    .m_axis_tkeep(remote_in_reg_m_axis_tkeep),
    .m_axis_tready(remote_in_reg_m_axis_tready),
    .m_axis_tlast(remote_in_reg_m_axis_tlast)
  );
  Arbiter switch_level1 ( // @[bfs_remote.scala 704:29]
    .io_in_0_ready(switch_level1_io_in_0_ready),
    .io_in_0_valid(switch_level1_io_in_0_valid),
    .io_in_0_bits_tdata(switch_level1_io_in_0_bits_tdata),
    .io_in_0_bits_tkeep(switch_level1_io_in_0_bits_tkeep),
    .io_in_0_bits_tlast(switch_level1_io_in_0_bits_tlast),
    .io_in_1_ready(switch_level1_io_in_1_ready),
    .io_in_1_valid(switch_level1_io_in_1_valid),
    .io_in_1_bits_tdata(switch_level1_io_in_1_bits_tdata),
    .io_in_1_bits_tkeep(switch_level1_io_in_1_bits_tkeep),
    .io_in_1_bits_tlast(switch_level1_io_in_1_bits_tlast),
    .io_out_ready(switch_level1_io_out_ready),
    .io_out_valid(switch_level1_io_out_valid),
    .io_out_bits_tdata(switch_level1_io_out_bits_tdata),
    .io_out_bits_tkeep(switch_level1_io_out_bits_tkeep),
    .io_out_bits_tlast(switch_level1_io_out_bits_tlast)
  );
  Remote_xbar_reg_slice mid ( // @[bfs_remote.scala 724:19]
    .aclk(mid_aclk),
    .aresetn(mid_aresetn),
    .s_axis_tdata(mid_s_axis_tdata),
    .s_axis_tvalid(mid_s_axis_tvalid),
    .s_axis_tkeep(mid_s_axis_tkeep),
    .s_axis_tready(mid_s_axis_tready),
    .s_axis_tlast(mid_s_axis_tlast),
    .m_axis_tdata(mid_m_axis_tdata),
    .m_axis_tvalid(mid_m_axis_tvalid),
    .m_axis_tkeep(mid_m_axis_tkeep),
    .m_axis_tready(mid_m_axis_tready),
    .m_axis_tlast(mid_m_axis_tlast)
  );
  axis_broadcaster_level1 xbar_level1 ( // @[bfs_remote.scala 733:27]
    .aclk(xbar_level1_aclk),
    .aresetn(xbar_level1_aresetn),
    .s_axis_tdata(xbar_level1_s_axis_tdata),
    .s_axis_tvalid(xbar_level1_s_axis_tvalid),
    .s_axis_tkeep(xbar_level1_s_axis_tkeep),
    .s_axis_tready(xbar_level1_s_axis_tready),
    .s_axis_tlast(xbar_level1_s_axis_tlast),
    .s_axis_tid(xbar_level1_s_axis_tid),
    .m_axis_tdata(xbar_level1_m_axis_tdata),
    .m_axis_tvalid(xbar_level1_m_axis_tvalid),
    .m_axis_tkeep(xbar_level1_m_axis_tkeep),
    .m_axis_tready(xbar_level1_m_axis_tready),
    .m_axis_tlast(xbar_level1_m_axis_tlast),
    .m_axis_tid(xbar_level1_m_axis_tid)
  );
  Remote_xbar_reg_slice backend_0 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_0_aclk),
    .aresetn(backend_0_aresetn),
    .s_axis_tdata(backend_0_s_axis_tdata),
    .s_axis_tvalid(backend_0_s_axis_tvalid),
    .s_axis_tkeep(backend_0_s_axis_tkeep),
    .s_axis_tready(backend_0_s_axis_tready),
    .s_axis_tlast(backend_0_s_axis_tlast),
    .m_axis_tdata(backend_0_m_axis_tdata),
    .m_axis_tvalid(backend_0_m_axis_tvalid),
    .m_axis_tkeep(backend_0_m_axis_tkeep),
    .m_axis_tready(backend_0_m_axis_tready),
    .m_axis_tlast(backend_0_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_1 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_1_aclk),
    .aresetn(backend_1_aresetn),
    .s_axis_tdata(backend_1_s_axis_tdata),
    .s_axis_tvalid(backend_1_s_axis_tvalid),
    .s_axis_tkeep(backend_1_s_axis_tkeep),
    .s_axis_tready(backend_1_s_axis_tready),
    .s_axis_tlast(backend_1_s_axis_tlast),
    .m_axis_tdata(backend_1_m_axis_tdata),
    .m_axis_tvalid(backend_1_m_axis_tvalid),
    .m_axis_tkeep(backend_1_m_axis_tkeep),
    .m_axis_tready(backend_1_m_axis_tready),
    .m_axis_tlast(backend_1_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_2 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_2_aclk),
    .aresetn(backend_2_aresetn),
    .s_axis_tdata(backend_2_s_axis_tdata),
    .s_axis_tvalid(backend_2_s_axis_tvalid),
    .s_axis_tkeep(backend_2_s_axis_tkeep),
    .s_axis_tready(backend_2_s_axis_tready),
    .s_axis_tlast(backend_2_s_axis_tlast),
    .m_axis_tdata(backend_2_m_axis_tdata),
    .m_axis_tvalid(backend_2_m_axis_tvalid),
    .m_axis_tkeep(backend_2_m_axis_tkeep),
    .m_axis_tready(backend_2_m_axis_tready),
    .m_axis_tlast(backend_2_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_3 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_3_aclk),
    .aresetn(backend_3_aresetn),
    .s_axis_tdata(backend_3_s_axis_tdata),
    .s_axis_tvalid(backend_3_s_axis_tvalid),
    .s_axis_tkeep(backend_3_s_axis_tkeep),
    .s_axis_tready(backend_3_s_axis_tready),
    .s_axis_tlast(backend_3_s_axis_tlast),
    .m_axis_tdata(backend_3_m_axis_tdata),
    .m_axis_tvalid(backend_3_m_axis_tvalid),
    .m_axis_tkeep(backend_3_m_axis_tkeep),
    .m_axis_tready(backend_3_m_axis_tready),
    .m_axis_tlast(backend_3_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_4 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_4_aclk),
    .aresetn(backend_4_aresetn),
    .s_axis_tdata(backend_4_s_axis_tdata),
    .s_axis_tvalid(backend_4_s_axis_tvalid),
    .s_axis_tkeep(backend_4_s_axis_tkeep),
    .s_axis_tready(backend_4_s_axis_tready),
    .s_axis_tlast(backend_4_s_axis_tlast),
    .m_axis_tdata(backend_4_m_axis_tdata),
    .m_axis_tvalid(backend_4_m_axis_tvalid),
    .m_axis_tkeep(backend_4_m_axis_tkeep),
    .m_axis_tready(backend_4_m_axis_tready),
    .m_axis_tlast(backend_4_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_5 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_5_aclk),
    .aresetn(backend_5_aresetn),
    .s_axis_tdata(backend_5_s_axis_tdata),
    .s_axis_tvalid(backend_5_s_axis_tvalid),
    .s_axis_tkeep(backend_5_s_axis_tkeep),
    .s_axis_tready(backend_5_s_axis_tready),
    .s_axis_tlast(backend_5_s_axis_tlast),
    .m_axis_tdata(backend_5_m_axis_tdata),
    .m_axis_tvalid(backend_5_m_axis_tvalid),
    .m_axis_tkeep(backend_5_m_axis_tkeep),
    .m_axis_tready(backend_5_m_axis_tready),
    .m_axis_tlast(backend_5_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_6 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_6_aclk),
    .aresetn(backend_6_aresetn),
    .s_axis_tdata(backend_6_s_axis_tdata),
    .s_axis_tvalid(backend_6_s_axis_tvalid),
    .s_axis_tkeep(backend_6_s_axis_tkeep),
    .s_axis_tready(backend_6_s_axis_tready),
    .s_axis_tlast(backend_6_s_axis_tlast),
    .m_axis_tdata(backend_6_m_axis_tdata),
    .m_axis_tvalid(backend_6_m_axis_tvalid),
    .m_axis_tkeep(backend_6_m_axis_tkeep),
    .m_axis_tready(backend_6_m_axis_tready),
    .m_axis_tlast(backend_6_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_7 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_7_aclk),
    .aresetn(backend_7_aresetn),
    .s_axis_tdata(backend_7_s_axis_tdata),
    .s_axis_tvalid(backend_7_s_axis_tvalid),
    .s_axis_tkeep(backend_7_s_axis_tkeep),
    .s_axis_tready(backend_7_s_axis_tready),
    .s_axis_tlast(backend_7_s_axis_tlast),
    .m_axis_tdata(backend_7_m_axis_tdata),
    .m_axis_tvalid(backend_7_m_axis_tvalid),
    .m_axis_tkeep(backend_7_m_axis_tkeep),
    .m_axis_tready(backend_7_m_axis_tready),
    .m_axis_tlast(backend_7_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_8 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_8_aclk),
    .aresetn(backend_8_aresetn),
    .s_axis_tdata(backend_8_s_axis_tdata),
    .s_axis_tvalid(backend_8_s_axis_tvalid),
    .s_axis_tkeep(backend_8_s_axis_tkeep),
    .s_axis_tready(backend_8_s_axis_tready),
    .s_axis_tlast(backend_8_s_axis_tlast),
    .m_axis_tdata(backend_8_m_axis_tdata),
    .m_axis_tvalid(backend_8_m_axis_tvalid),
    .m_axis_tkeep(backend_8_m_axis_tkeep),
    .m_axis_tready(backend_8_m_axis_tready),
    .m_axis_tlast(backend_8_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_9 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_9_aclk),
    .aresetn(backend_9_aresetn),
    .s_axis_tdata(backend_9_s_axis_tdata),
    .s_axis_tvalid(backend_9_s_axis_tvalid),
    .s_axis_tkeep(backend_9_s_axis_tkeep),
    .s_axis_tready(backend_9_s_axis_tready),
    .s_axis_tlast(backend_9_s_axis_tlast),
    .m_axis_tdata(backend_9_m_axis_tdata),
    .m_axis_tvalid(backend_9_m_axis_tvalid),
    .m_axis_tkeep(backend_9_m_axis_tkeep),
    .m_axis_tready(backend_9_m_axis_tready),
    .m_axis_tlast(backend_9_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_10 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_10_aclk),
    .aresetn(backend_10_aresetn),
    .s_axis_tdata(backend_10_s_axis_tdata),
    .s_axis_tvalid(backend_10_s_axis_tvalid),
    .s_axis_tkeep(backend_10_s_axis_tkeep),
    .s_axis_tready(backend_10_s_axis_tready),
    .s_axis_tlast(backend_10_s_axis_tlast),
    .m_axis_tdata(backend_10_m_axis_tdata),
    .m_axis_tvalid(backend_10_m_axis_tvalid),
    .m_axis_tkeep(backend_10_m_axis_tkeep),
    .m_axis_tready(backend_10_m_axis_tready),
    .m_axis_tlast(backend_10_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_11 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_11_aclk),
    .aresetn(backend_11_aresetn),
    .s_axis_tdata(backend_11_s_axis_tdata),
    .s_axis_tvalid(backend_11_s_axis_tvalid),
    .s_axis_tkeep(backend_11_s_axis_tkeep),
    .s_axis_tready(backend_11_s_axis_tready),
    .s_axis_tlast(backend_11_s_axis_tlast),
    .m_axis_tdata(backend_11_m_axis_tdata),
    .m_axis_tvalid(backend_11_m_axis_tvalid),
    .m_axis_tkeep(backend_11_m_axis_tkeep),
    .m_axis_tready(backend_11_m_axis_tready),
    .m_axis_tlast(backend_11_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_12 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_12_aclk),
    .aresetn(backend_12_aresetn),
    .s_axis_tdata(backend_12_s_axis_tdata),
    .s_axis_tvalid(backend_12_s_axis_tvalid),
    .s_axis_tkeep(backend_12_s_axis_tkeep),
    .s_axis_tready(backend_12_s_axis_tready),
    .s_axis_tlast(backend_12_s_axis_tlast),
    .m_axis_tdata(backend_12_m_axis_tdata),
    .m_axis_tvalid(backend_12_m_axis_tvalid),
    .m_axis_tkeep(backend_12_m_axis_tkeep),
    .m_axis_tready(backend_12_m_axis_tready),
    .m_axis_tlast(backend_12_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_13 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_13_aclk),
    .aresetn(backend_13_aresetn),
    .s_axis_tdata(backend_13_s_axis_tdata),
    .s_axis_tvalid(backend_13_s_axis_tvalid),
    .s_axis_tkeep(backend_13_s_axis_tkeep),
    .s_axis_tready(backend_13_s_axis_tready),
    .s_axis_tlast(backend_13_s_axis_tlast),
    .m_axis_tdata(backend_13_m_axis_tdata),
    .m_axis_tvalid(backend_13_m_axis_tvalid),
    .m_axis_tkeep(backend_13_m_axis_tkeep),
    .m_axis_tready(backend_13_m_axis_tready),
    .m_axis_tlast(backend_13_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_14 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_14_aclk),
    .aresetn(backend_14_aresetn),
    .s_axis_tdata(backend_14_s_axis_tdata),
    .s_axis_tvalid(backend_14_s_axis_tvalid),
    .s_axis_tkeep(backend_14_s_axis_tkeep),
    .s_axis_tready(backend_14_s_axis_tready),
    .s_axis_tlast(backend_14_s_axis_tlast),
    .m_axis_tdata(backend_14_m_axis_tdata),
    .m_axis_tvalid(backend_14_m_axis_tvalid),
    .m_axis_tkeep(backend_14_m_axis_tkeep),
    .m_axis_tready(backend_14_m_axis_tready),
    .m_axis_tlast(backend_14_m_axis_tlast)
  );
  Remote_xbar_reg_slice backend_15 ( // @[bfs_remote.scala 741:43]
    .aclk(backend_15_aclk),
    .aresetn(backend_15_aresetn),
    .s_axis_tdata(backend_15_s_axis_tdata),
    .s_axis_tvalid(backend_15_s_axis_tvalid),
    .s_axis_tkeep(backend_15_s_axis_tkeep),
    .s_axis_tready(backend_15_s_axis_tready),
    .s_axis_tlast(backend_15_s_axis_tlast),
    .m_axis_tdata(backend_15_m_axis_tdata),
    .m_axis_tvalid(backend_15_m_axis_tvalid),
    .m_axis_tkeep(backend_15_m_axis_tkeep),
    .m_axis_tready(backend_15_m_axis_tready),
    .m_axis_tlast(backend_15_m_axis_tlast)
  );
  assign io_ddr_in_0_ready = combiner_level0_s_axis_tready[0]; // @[bfs_remote.scala 637:65]
  assign io_ddr_in_1_ready = combiner_level0_s_axis_tready[1]; // @[bfs_remote.scala 637:65]
  assign io_ddr_in_2_ready = combiner_level0_s_axis_tready[2]; // @[bfs_remote.scala 637:65]
  assign io_ddr_in_3_ready = combiner_level0_s_axis_tready[3]; // @[bfs_remote.scala 637:65]
  assign io_pe_out_0_valid = backend_0_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_0_bits_tdata = backend_0_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_0_bits_tkeep = _io_pe_out_0_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_0_bits_tlast = backend_0_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_1_valid = backend_1_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_1_bits_tdata = backend_1_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_1_bits_tkeep = _io_pe_out_1_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_1_bits_tlast = backend_1_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_2_valid = backend_2_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_2_bits_tdata = backend_2_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_2_bits_tkeep = _io_pe_out_2_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_2_bits_tlast = backend_2_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_3_valid = backend_3_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_3_bits_tdata = backend_3_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_3_bits_tkeep = _io_pe_out_3_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_3_bits_tlast = backend_3_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_4_valid = backend_4_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_4_bits_tdata = backend_4_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_4_bits_tkeep = _io_pe_out_4_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_4_bits_tlast = backend_4_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_5_valid = backend_5_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_5_bits_tdata = backend_5_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_5_bits_tkeep = _io_pe_out_5_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_5_bits_tlast = backend_5_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_6_valid = backend_6_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_6_bits_tdata = backend_6_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_6_bits_tkeep = _io_pe_out_6_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_6_bits_tlast = backend_6_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_7_valid = backend_7_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_7_bits_tdata = backend_7_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_7_bits_tkeep = _io_pe_out_7_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_7_bits_tlast = backend_7_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_8_valid = backend_8_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_8_bits_tdata = backend_8_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_8_bits_tkeep = _io_pe_out_8_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_8_bits_tlast = backend_8_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_9_valid = backend_9_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_9_bits_tdata = backend_9_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_9_bits_tkeep = _io_pe_out_9_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_9_bits_tlast = backend_9_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_10_valid = backend_10_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_10_bits_tdata = backend_10_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_10_bits_tkeep = _io_pe_out_10_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_10_bits_tlast = backend_10_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_11_valid = backend_11_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_11_bits_tdata = backend_11_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_11_bits_tkeep = _io_pe_out_11_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_11_bits_tlast = backend_11_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_12_valid = backend_12_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_12_bits_tdata = backend_12_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_12_bits_tkeep = _io_pe_out_12_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_12_bits_tlast = backend_12_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_13_valid = backend_13_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_13_bits_tdata = backend_13_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_13_bits_tkeep = _io_pe_out_13_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_13_bits_tlast = backend_13_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_14_valid = backend_14_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_14_bits_tdata = backend_14_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_14_bits_tkeep = _io_pe_out_14_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_14_bits_tlast = backend_14_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_pe_out_15_valid = backend_15_m_axis_tvalid; // @[bfs_remote.scala 758:16]
  assign io_pe_out_15_bits_tdata = backend_15_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign io_pe_out_15_bits_tkeep = _io_pe_out_15_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 127:13]
  assign io_pe_out_15_bits_tlast = backend_15_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign io_remote_out_0_valid = xbar_level0_m_axis_tvalid[1]; // @[bfs_remote.scala 659:46]
  assign io_remote_out_0_bits_tdata = xbar_level0_m_axis_tdata[1023:512]; // @[nf_arm_doce_top.scala 125:21]
  assign io_remote_out_0_bits_tkeep = xbar_level0_m_axis_tkeep[79:64]; // @[nf_arm_doce_top.scala 127:13]
  assign io_remote_out_1_valid = xbar_level0_m_axis_tvalid[2]; // @[bfs_remote.scala 659:46]
  assign io_remote_out_1_bits_tdata = xbar_level0_m_axis_tdata[1535:1024]; // @[nf_arm_doce_top.scala 125:21]
  assign io_remote_out_1_bits_tkeep = xbar_level0_m_axis_tkeep[143:128]; // @[nf_arm_doce_top.scala 127:13]
  assign io_remote_out_2_valid = xbar_level0_m_axis_tvalid[3]; // @[bfs_remote.scala 659:46]
  assign io_remote_out_2_bits_tdata = xbar_level0_m_axis_tdata[2047:1536]; // @[nf_arm_doce_top.scala 125:21]
  assign io_remote_out_2_bits_tkeep = xbar_level0_m_axis_tkeep[207:192]; // @[nf_arm_doce_top.scala 127:13]
  assign io_remote_out_3_valid = xbar_level0_m_axis_tvalid[4]; // @[bfs_remote.scala 659:46]
  assign io_remote_out_3_bits_tdata = xbar_level0_m_axis_tdata[2559:2048]; // @[nf_arm_doce_top.scala 125:21]
  assign io_remote_out_3_bits_tkeep = xbar_level0_m_axis_tkeep[271:256]; // @[nf_arm_doce_top.scala 127:13]
  assign io_remote_in_ready = remote_in_reg_s_axis_tready; // @[bfs_remote.scala 701:22]
  assign combiner_level0_aclk = clock; // @[bfs_remote.scala 629:42]
  assign combiner_level0_aresetn = ~reset; // @[bfs_remote.scala 630:33]
  assign combiner_level0_s_axis_tdata = {combiner_level0_io_s_axis_tdata_hi,combiner_level0_io_s_axis_tdata_lo}; // @[bfs_remote.scala 631:103]
  assign combiner_level0_s_axis_tvalid = {combiner_level0_io_s_axis_tvalid_lo,combiner_level0_io_s_axis_tvalid_lo}; // @[bfs_remote.scala 635:116]
  assign combiner_level0_s_axis_tkeep = {{48'd0}, _combiner_level0_io_s_axis_tkeep_T_32}; // @[bfs_remote.scala 633:33]
  assign combiner_level0_s_axis_tlast = {combiner_level0_io_s_axis_tlast_hi,combiner_level0_io_s_axis_tlast_lo}; // @[bfs_remote.scala 634:103]
  assign combiner_level0_s_axis_tid = 4'h0;
  assign combiner_level0_m_axis_tready = frontend_s_axis_tready; // @[bfs_remote.scala 647:36]
  assign frontend_aclk = clock; // @[bfs_remote.scala 641:35]
  assign frontend_aresetn = ~reset; // @[bfs_remote.scala 642:26]
  assign frontend_s_axis_tdata = combiner_level0_m_axis_tdata; // @[bfs_remote.scala 644:28]
  assign frontend_s_axis_tvalid = combiner_level0_m_axis_tvalid; // @[bfs_remote.scala 643:29]
  assign frontend_s_axis_tkeep = combiner_level0_m_axis_tkeep; // @[bfs_remote.scala 645:28]
  assign frontend_s_axis_tlast = combiner_level0_m_axis_tlast; // @[bfs_remote.scala 646:28]
  assign frontend_m_axis_tready = xbar_level0_s_axis_tready; // @[bfs_remote.scala 655:29]
  assign xbar_level0_aclk = clock; // @[bfs_remote.scala 650:38]
  assign xbar_level0_aresetn = ~reset; // @[bfs_remote.scala 651:29]
  assign xbar_level0_s_axis_tdata = frontend_m_axis_tdata; // @[bfs_remote.scala 652:31]
  assign xbar_level0_s_axis_tvalid = frontend_m_axis_tvalid; // @[bfs_remote.scala 653:32]
  assign xbar_level0_s_axis_tkeep = {xbar_level0_io_s_axis_tkeep_hi,xbar_level0_io_s_axis_tkeep_lo}; // @[bfs_remote.scala 654:124]
  assign xbar_level0_s_axis_tlast = 1'h0;
  assign xbar_level0_s_axis_tid = 1'h0;
  assign xbar_level0_m_axis_tready = {xbar_level0_io_m_axis_tready_hi_1,collector_io_in_ready}; // @[Cat.scala 30:58]
  assign collector_clock = clock;
  assign collector_reset = reset;
  assign collector_io_in_valid = xbar_level0_m_axis_tvalid[0]; // @[bfs_remote.scala 683:56]
  assign collector_io_in_bits_tdata = xbar_level0_m_axis_tdata[511:0]; // @[bfs_remote.scala 685:60]
  assign collector_io_in_bits_tkeep = {collector_io_in_bits_tkeep_hi,collector_io_in_bits_tkeep_lo}; // @[bfs_remote.scala 684:53]
  assign collector_io_out_ready = buffer1_s_axis_tready; // @[bfs_remote.scala 695:26]
  assign collector_io_flush = flush_reg; // @[bfs_remote.scala 688:22]
  assign buffer1_s_axis_aclk = clock; // @[bfs_remote.scala 691:41]
  assign buffer1_s_axis_aresetn = ~reset; // @[bfs_remote.scala 692:32]
  assign buffer1_s_axis_tdata = collector_io_out_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign buffer1_s_axis_tvalid = collector_io_out_valid; // @[bfs_remote.scala 694:28]
  assign buffer1_s_axis_tkeep = {{48'd0}, collector_io_out_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign buffer1_s_axis_tlast = collector_io_out_bits_tlast; // @[nf_arm_doce_top.scala 120:11]
  assign buffer1_s_axis_tid = 1'h0;
  assign buffer1_m_axis_tready = switch_level1_io_in_1_ready; // @[bfs_remote.scala 707:28]
  assign remote_in_reg_aclk = clock; // @[bfs_remote.scala 698:40]
  assign remote_in_reg_aresetn = ~reset; // @[bfs_remote.scala 699:31]
  assign remote_in_reg_s_axis_tdata = io_remote_in_bits_tdata; // @[nf_arm_doce_top.scala 119:11]
  assign remote_in_reg_s_axis_tvalid = io_remote_in_valid; // @[bfs_remote.scala 702:34]
  assign remote_in_reg_s_axis_tkeep = {{48'd0}, io_remote_in_bits_tkeep}; // @[nf_arm_doce_top.scala 121:11]
  assign remote_in_reg_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 120:11]
  assign remote_in_reg_m_axis_tready = switch_level1_io_in_0_ready; // @[bfs_remote.scala 710:34]
  assign switch_level1_io_in_0_valid = remote_in_reg_m_axis_tvalid; // @[bfs_remote.scala 709:32]
  assign switch_level1_io_in_0_bits_tdata = remote_in_reg_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign switch_level1_io_in_0_bits_tkeep = remote_in_reg_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  assign switch_level1_io_in_0_bits_tlast = remote_in_reg_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign switch_level1_io_in_1_valid = buffer1_m_axis_tvalid; // @[bfs_remote.scala 706:32]
  assign switch_level1_io_in_1_bits_tdata = buffer1_m_axis_tdata; // @[nf_arm_doce_top.scala 125:21]
  assign switch_level1_io_in_1_bits_tkeep = buffer1_m_axis_tkeep; // @[nf_arm_doce_top.scala 127:21]
  assign switch_level1_io_in_1_bits_tlast = buffer1_m_axis_tlast; // @[nf_arm_doce_top.scala 126:21]
  assign switch_level1_io_out_ready = mid_s_axis_tready; // @[bfs_remote.scala 731:30]
  assign mid_aclk = clock; // @[bfs_remote.scala 725:30]
  assign mid_aresetn = ~reset; // @[bfs_remote.scala 726:21]
  assign mid_s_axis_tdata = switch_level1_io_out_bits_tdata; // @[bfs_remote.scala 728:23]
  assign mid_s_axis_tvalid = switch_level1_io_out_valid; // @[bfs_remote.scala 727:24]
  assign mid_s_axis_tkeep = switch_level1_io_out_bits_tkeep & _GEN_2; // @[bfs_remote.scala 730:58]
  assign mid_s_axis_tlast = switch_level1_io_out_bits_tlast; // @[bfs_remote.scala 729:23]
  assign mid_m_axis_tready = xbar_level1_s_axis_tready; // @[bfs_remote.scala 739:24]
  assign xbar_level1_aclk = clock; // @[bfs_remote.scala 734:38]
  assign xbar_level1_aresetn = ~reset; // @[bfs_remote.scala 735:29]
  assign xbar_level1_s_axis_tdata = mid_m_axis_tdata; // @[bfs_remote.scala 736:31]
  assign xbar_level1_s_axis_tvalid = mid_m_axis_tvalid; // @[bfs_remote.scala 737:32]
  assign xbar_level1_s_axis_tkeep = {xbar_level1_io_s_axis_tkeep_hi,xbar_level1_io_s_axis_tkeep_lo}; // @[bfs_remote.scala 738:114]
  assign xbar_level1_s_axis_tlast = 1'h0;
  assign xbar_level1_s_axis_tid = 1'h0;
  assign xbar_level1_m_axis_tready = {xbar_level1_io_m_axis_tready_hi,xbar_level1_io_m_axis_tready_lo}; // @[bfs_remote.scala 754:12]
  assign backend_0_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_0_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_0_s_axis_tdata = xbar_level1_m_axis_tdata[511:0]; // @[bfs_remote.scala 746:55]
  assign backend_0_s_axis_tvalid = xbar_level1_m_axis_tvalid[0]; // @[bfs_remote.scala 749:57]
  assign backend_0_s_axis_tkeep = xbar_level1_m_axis_tkeep[63:0]; // @[bfs_remote.scala 747:55]
  assign backend_0_s_axis_tlast = xbar_level1_m_axis_tlast[0]; // @[bfs_remote.scala 748:55]
  assign backend_0_m_axis_tready = io_pe_out_0_ready; // @[bfs_remote.scala 759:35]
  assign backend_1_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_1_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_1_s_axis_tdata = xbar_level1_m_axis_tdata[1023:512]; // @[bfs_remote.scala 746:55]
  assign backend_1_s_axis_tvalid = xbar_level1_m_axis_tvalid[1]; // @[bfs_remote.scala 749:57]
  assign backend_1_s_axis_tkeep = xbar_level1_m_axis_tkeep[127:64]; // @[bfs_remote.scala 747:55]
  assign backend_1_s_axis_tlast = xbar_level1_m_axis_tlast[1]; // @[bfs_remote.scala 748:55]
  assign backend_1_m_axis_tready = io_pe_out_1_ready; // @[bfs_remote.scala 759:35]
  assign backend_2_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_2_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_2_s_axis_tdata = xbar_level1_m_axis_tdata[1535:1024]; // @[bfs_remote.scala 746:55]
  assign backend_2_s_axis_tvalid = xbar_level1_m_axis_tvalid[2]; // @[bfs_remote.scala 749:57]
  assign backend_2_s_axis_tkeep = xbar_level1_m_axis_tkeep[191:128]; // @[bfs_remote.scala 747:55]
  assign backend_2_s_axis_tlast = xbar_level1_m_axis_tlast[2]; // @[bfs_remote.scala 748:55]
  assign backend_2_m_axis_tready = io_pe_out_2_ready; // @[bfs_remote.scala 759:35]
  assign backend_3_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_3_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_3_s_axis_tdata = xbar_level1_m_axis_tdata[2047:1536]; // @[bfs_remote.scala 746:55]
  assign backend_3_s_axis_tvalid = xbar_level1_m_axis_tvalid[3]; // @[bfs_remote.scala 749:57]
  assign backend_3_s_axis_tkeep = xbar_level1_m_axis_tkeep[255:192]; // @[bfs_remote.scala 747:55]
  assign backend_3_s_axis_tlast = xbar_level1_m_axis_tlast[3]; // @[bfs_remote.scala 748:55]
  assign backend_3_m_axis_tready = io_pe_out_3_ready; // @[bfs_remote.scala 759:35]
  assign backend_4_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_4_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_4_s_axis_tdata = xbar_level1_m_axis_tdata[2559:2048]; // @[bfs_remote.scala 746:55]
  assign backend_4_s_axis_tvalid = xbar_level1_m_axis_tvalid[4]; // @[bfs_remote.scala 749:57]
  assign backend_4_s_axis_tkeep = xbar_level1_m_axis_tkeep[319:256]; // @[bfs_remote.scala 747:55]
  assign backend_4_s_axis_tlast = xbar_level1_m_axis_tlast[4]; // @[bfs_remote.scala 748:55]
  assign backend_4_m_axis_tready = io_pe_out_4_ready; // @[bfs_remote.scala 759:35]
  assign backend_5_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_5_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_5_s_axis_tdata = xbar_level1_m_axis_tdata[3071:2560]; // @[bfs_remote.scala 746:55]
  assign backend_5_s_axis_tvalid = xbar_level1_m_axis_tvalid[5]; // @[bfs_remote.scala 749:57]
  assign backend_5_s_axis_tkeep = xbar_level1_m_axis_tkeep[383:320]; // @[bfs_remote.scala 747:55]
  assign backend_5_s_axis_tlast = xbar_level1_m_axis_tlast[5]; // @[bfs_remote.scala 748:55]
  assign backend_5_m_axis_tready = io_pe_out_5_ready; // @[bfs_remote.scala 759:35]
  assign backend_6_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_6_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_6_s_axis_tdata = xbar_level1_m_axis_tdata[3583:3072]; // @[bfs_remote.scala 746:55]
  assign backend_6_s_axis_tvalid = xbar_level1_m_axis_tvalid[6]; // @[bfs_remote.scala 749:57]
  assign backend_6_s_axis_tkeep = xbar_level1_m_axis_tkeep[447:384]; // @[bfs_remote.scala 747:55]
  assign backend_6_s_axis_tlast = xbar_level1_m_axis_tlast[6]; // @[bfs_remote.scala 748:55]
  assign backend_6_m_axis_tready = io_pe_out_6_ready; // @[bfs_remote.scala 759:35]
  assign backend_7_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_7_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_7_s_axis_tdata = xbar_level1_m_axis_tdata[4095:3584]; // @[bfs_remote.scala 746:55]
  assign backend_7_s_axis_tvalid = xbar_level1_m_axis_tvalid[7]; // @[bfs_remote.scala 749:57]
  assign backend_7_s_axis_tkeep = xbar_level1_m_axis_tkeep[511:448]; // @[bfs_remote.scala 747:55]
  assign backend_7_s_axis_tlast = xbar_level1_m_axis_tlast[7]; // @[bfs_remote.scala 748:55]
  assign backend_7_m_axis_tready = io_pe_out_7_ready; // @[bfs_remote.scala 759:35]
  assign backend_8_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_8_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_8_s_axis_tdata = xbar_level1_m_axis_tdata[4607:4096]; // @[bfs_remote.scala 746:55]
  assign backend_8_s_axis_tvalid = xbar_level1_m_axis_tvalid[8]; // @[bfs_remote.scala 749:57]
  assign backend_8_s_axis_tkeep = xbar_level1_m_axis_tkeep[575:512]; // @[bfs_remote.scala 747:55]
  assign backend_8_s_axis_tlast = xbar_level1_m_axis_tlast[8]; // @[bfs_remote.scala 748:55]
  assign backend_8_m_axis_tready = io_pe_out_8_ready; // @[bfs_remote.scala 759:35]
  assign backend_9_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_9_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_9_s_axis_tdata = xbar_level1_m_axis_tdata[5119:4608]; // @[bfs_remote.scala 746:55]
  assign backend_9_s_axis_tvalid = xbar_level1_m_axis_tvalid[9]; // @[bfs_remote.scala 749:57]
  assign backend_9_s_axis_tkeep = xbar_level1_m_axis_tkeep[639:576]; // @[bfs_remote.scala 747:55]
  assign backend_9_s_axis_tlast = xbar_level1_m_axis_tlast[9]; // @[bfs_remote.scala 748:55]
  assign backend_9_m_axis_tready = io_pe_out_9_ready; // @[bfs_remote.scala 759:35]
  assign backend_10_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_10_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_10_s_axis_tdata = xbar_level1_m_axis_tdata[5631:5120]; // @[bfs_remote.scala 746:55]
  assign backend_10_s_axis_tvalid = xbar_level1_m_axis_tvalid[10]; // @[bfs_remote.scala 749:57]
  assign backend_10_s_axis_tkeep = xbar_level1_m_axis_tkeep[703:640]; // @[bfs_remote.scala 747:55]
  assign backend_10_s_axis_tlast = xbar_level1_m_axis_tlast[10]; // @[bfs_remote.scala 748:55]
  assign backend_10_m_axis_tready = io_pe_out_10_ready; // @[bfs_remote.scala 759:35]
  assign backend_11_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_11_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_11_s_axis_tdata = xbar_level1_m_axis_tdata[6143:5632]; // @[bfs_remote.scala 746:55]
  assign backend_11_s_axis_tvalid = xbar_level1_m_axis_tvalid[11]; // @[bfs_remote.scala 749:57]
  assign backend_11_s_axis_tkeep = xbar_level1_m_axis_tkeep[767:704]; // @[bfs_remote.scala 747:55]
  assign backend_11_s_axis_tlast = xbar_level1_m_axis_tlast[11]; // @[bfs_remote.scala 748:55]
  assign backend_11_m_axis_tready = io_pe_out_11_ready; // @[bfs_remote.scala 759:35]
  assign backend_12_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_12_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_12_s_axis_tdata = xbar_level1_m_axis_tdata[6655:6144]; // @[bfs_remote.scala 746:55]
  assign backend_12_s_axis_tvalid = xbar_level1_m_axis_tvalid[12]; // @[bfs_remote.scala 749:57]
  assign backend_12_s_axis_tkeep = xbar_level1_m_axis_tkeep[831:768]; // @[bfs_remote.scala 747:55]
  assign backend_12_s_axis_tlast = xbar_level1_m_axis_tlast[12]; // @[bfs_remote.scala 748:55]
  assign backend_12_m_axis_tready = io_pe_out_12_ready; // @[bfs_remote.scala 759:35]
  assign backend_13_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_13_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_13_s_axis_tdata = xbar_level1_m_axis_tdata[7167:6656]; // @[bfs_remote.scala 746:55]
  assign backend_13_s_axis_tvalid = xbar_level1_m_axis_tvalid[13]; // @[bfs_remote.scala 749:57]
  assign backend_13_s_axis_tkeep = xbar_level1_m_axis_tkeep[895:832]; // @[bfs_remote.scala 747:55]
  assign backend_13_s_axis_tlast = xbar_level1_m_axis_tlast[13]; // @[bfs_remote.scala 748:55]
  assign backend_13_m_axis_tready = io_pe_out_13_ready; // @[bfs_remote.scala 759:35]
  assign backend_14_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_14_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_14_s_axis_tdata = xbar_level1_m_axis_tdata[7679:7168]; // @[bfs_remote.scala 746:55]
  assign backend_14_s_axis_tvalid = xbar_level1_m_axis_tvalid[14]; // @[bfs_remote.scala 749:57]
  assign backend_14_s_axis_tkeep = xbar_level1_m_axis_tkeep[959:896]; // @[bfs_remote.scala 747:55]
  assign backend_14_s_axis_tlast = xbar_level1_m_axis_tlast[14]; // @[bfs_remote.scala 748:55]
  assign backend_14_m_axis_tready = io_pe_out_14_ready; // @[bfs_remote.scala 759:35]
  assign backend_15_aclk = clock; // @[bfs_remote.scala 744:32]
  assign backend_15_aresetn = ~reset; // @[bfs_remote.scala 745:23]
  assign backend_15_s_axis_tdata = xbar_level1_m_axis_tdata[8191:7680]; // @[bfs_remote.scala 746:55]
  assign backend_15_s_axis_tvalid = xbar_level1_m_axis_tvalid[15]; // @[bfs_remote.scala 749:57]
  assign backend_15_s_axis_tkeep = xbar_level1_m_axis_tkeep[1023:960]; // @[bfs_remote.scala 747:55]
  assign backend_15_s_axis_tlast = xbar_level1_m_axis_tlast[15]; // @[bfs_remote.scala 748:55]
  assign backend_15_m_axis_tready = io_pe_out_15_ready; // @[bfs_remote.scala 759:35]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 625:30]
      local_fpga_id <= 2'h0; // @[bfs_remote.scala 625:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[bfs_remote.scala 626:17]
    end
    if (reset) begin // @[bfs_remote.scala 676:26]
      flush_reg <= 1'h0; // @[bfs_remote.scala 676:26]
    end else if (io_signal) begin // @[bfs_remote.scala 677:18]
      flush_reg <= 1'h0; // @[bfs_remote.scala 678:15]
    end else begin
      flush_reg <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  flush_reg = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module flow_control(
  input          clock,
  input          reset,
  input  [511:0] io_data,
  input  [15:0]  io_keep,
  input          io_handshake,
  input          io_handshake_last,
  input  [31:0]  io_period,
  output         io_pending_valid,
  output [31:0]  io_pending_bits,
  input  [31:0]  io_parameter,
  input  [1:0]   io_idol_fpga_num
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  layer1_0_aclk; // @[bfs_remote.scala 208:34]
  wire  layer1_0_aresetn; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_0_s_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_0_s_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_0_s_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_0_s_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_0_s_axis_tlast; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_0_m_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_0_m_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_0_m_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_0_m_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_0_m_axis_tlast; // @[bfs_remote.scala 208:34]
  wire  layer1_1_aclk; // @[bfs_remote.scala 208:34]
  wire  layer1_1_aresetn; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_1_s_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_1_s_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_1_s_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_1_s_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_1_s_axis_tlast; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_1_m_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_1_m_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_1_m_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_1_m_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_1_m_axis_tlast; // @[bfs_remote.scala 208:34]
  wire  layer1_2_aclk; // @[bfs_remote.scala 208:34]
  wire  layer1_2_aresetn; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_2_s_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_2_s_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_2_s_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_2_s_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_2_s_axis_tlast; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_2_m_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_2_m_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_2_m_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_2_m_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_2_m_axis_tlast; // @[bfs_remote.scala 208:34]
  wire  layer1_3_aclk; // @[bfs_remote.scala 208:34]
  wire  layer1_3_aresetn; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_3_s_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_3_s_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_3_s_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_3_s_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_3_s_axis_tlast; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_3_m_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_3_m_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_3_m_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_3_m_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_3_m_axis_tlast; // @[bfs_remote.scala 208:34]
  wire  layer1_4_aclk; // @[bfs_remote.scala 208:34]
  wire  layer1_4_aresetn; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_4_s_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_4_s_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_4_s_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_4_s_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_4_s_axis_tlast; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_4_m_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_4_m_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_4_m_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_4_m_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_4_m_axis_tlast; // @[bfs_remote.scala 208:34]
  wire  layer1_5_aclk; // @[bfs_remote.scala 208:34]
  wire  layer1_5_aresetn; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_5_s_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_5_s_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_5_s_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_5_s_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_5_s_axis_tlast; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_5_m_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_5_m_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_5_m_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_5_m_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_5_m_axis_tlast; // @[bfs_remote.scala 208:34]
  wire  layer1_6_aclk; // @[bfs_remote.scala 208:34]
  wire  layer1_6_aresetn; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_6_s_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_6_s_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_6_s_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_6_s_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_6_s_axis_tlast; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_6_m_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_6_m_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_6_m_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_6_m_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_6_m_axis_tlast; // @[bfs_remote.scala 208:34]
  wire  layer1_7_aclk; // @[bfs_remote.scala 208:34]
  wire  layer1_7_aresetn; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_7_s_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_7_s_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_7_s_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_7_s_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_7_s_axis_tlast; // @[bfs_remote.scala 208:34]
  wire [31:0] layer1_7_m_axis_tdata; // @[bfs_remote.scala 208:34]
  wire  layer1_7_m_axis_tvalid; // @[bfs_remote.scala 208:34]
  wire [3:0] layer1_7_m_axis_tkeep; // @[bfs_remote.scala 208:34]
  wire  layer1_7_m_axis_tready; // @[bfs_remote.scala 208:34]
  wire  layer1_7_m_axis_tlast; // @[bfs_remote.scala 208:34]
  wire  layer2_0_aclk; // @[bfs_remote.scala 217:34]
  wire  layer2_0_aresetn; // @[bfs_remote.scala 217:34]
  wire [31:0] layer2_0_s_axis_tdata; // @[bfs_remote.scala 217:34]
  wire  layer2_0_s_axis_tvalid; // @[bfs_remote.scala 217:34]
  wire [3:0] layer2_0_s_axis_tkeep; // @[bfs_remote.scala 217:34]
  wire  layer2_0_s_axis_tready; // @[bfs_remote.scala 217:34]
  wire  layer2_0_s_axis_tlast; // @[bfs_remote.scala 217:34]
  wire [31:0] layer2_0_m_axis_tdata; // @[bfs_remote.scala 217:34]
  wire  layer2_0_m_axis_tvalid; // @[bfs_remote.scala 217:34]
  wire [3:0] layer2_0_m_axis_tkeep; // @[bfs_remote.scala 217:34]
  wire  layer2_0_m_axis_tready; // @[bfs_remote.scala 217:34]
  wire  layer2_0_m_axis_tlast; // @[bfs_remote.scala 217:34]
  wire  layer2_1_aclk; // @[bfs_remote.scala 217:34]
  wire  layer2_1_aresetn; // @[bfs_remote.scala 217:34]
  wire [31:0] layer2_1_s_axis_tdata; // @[bfs_remote.scala 217:34]
  wire  layer2_1_s_axis_tvalid; // @[bfs_remote.scala 217:34]
  wire [3:0] layer2_1_s_axis_tkeep; // @[bfs_remote.scala 217:34]
  wire  layer2_1_s_axis_tready; // @[bfs_remote.scala 217:34]
  wire  layer2_1_s_axis_tlast; // @[bfs_remote.scala 217:34]
  wire [31:0] layer2_1_m_axis_tdata; // @[bfs_remote.scala 217:34]
  wire  layer2_1_m_axis_tvalid; // @[bfs_remote.scala 217:34]
  wire [3:0] layer2_1_m_axis_tkeep; // @[bfs_remote.scala 217:34]
  wire  layer2_1_m_axis_tready; // @[bfs_remote.scala 217:34]
  wire  layer2_1_m_axis_tlast; // @[bfs_remote.scala 217:34]
  wire  layer2_2_aclk; // @[bfs_remote.scala 217:34]
  wire  layer2_2_aresetn; // @[bfs_remote.scala 217:34]
  wire [31:0] layer2_2_s_axis_tdata; // @[bfs_remote.scala 217:34]
  wire  layer2_2_s_axis_tvalid; // @[bfs_remote.scala 217:34]
  wire [3:0] layer2_2_s_axis_tkeep; // @[bfs_remote.scala 217:34]
  wire  layer2_2_s_axis_tready; // @[bfs_remote.scala 217:34]
  wire  layer2_2_s_axis_tlast; // @[bfs_remote.scala 217:34]
  wire [31:0] layer2_2_m_axis_tdata; // @[bfs_remote.scala 217:34]
  wire  layer2_2_m_axis_tvalid; // @[bfs_remote.scala 217:34]
  wire [3:0] layer2_2_m_axis_tkeep; // @[bfs_remote.scala 217:34]
  wire  layer2_2_m_axis_tready; // @[bfs_remote.scala 217:34]
  wire  layer2_2_m_axis_tlast; // @[bfs_remote.scala 217:34]
  wire  layer2_3_aclk; // @[bfs_remote.scala 217:34]
  wire  layer2_3_aresetn; // @[bfs_remote.scala 217:34]
  wire [31:0] layer2_3_s_axis_tdata; // @[bfs_remote.scala 217:34]
  wire  layer2_3_s_axis_tvalid; // @[bfs_remote.scala 217:34]
  wire [3:0] layer2_3_s_axis_tkeep; // @[bfs_remote.scala 217:34]
  wire  layer2_3_s_axis_tready; // @[bfs_remote.scala 217:34]
  wire  layer2_3_s_axis_tlast; // @[bfs_remote.scala 217:34]
  wire [31:0] layer2_3_m_axis_tdata; // @[bfs_remote.scala 217:34]
  wire  layer2_3_m_axis_tvalid; // @[bfs_remote.scala 217:34]
  wire [3:0] layer2_3_m_axis_tkeep; // @[bfs_remote.scala 217:34]
  wire  layer2_3_m_axis_tready; // @[bfs_remote.scala 217:34]
  wire  layer2_3_m_axis_tlast; // @[bfs_remote.scala 217:34]
  wire  layer3_0_aclk; // @[bfs_remote.scala 229:34]
  wire  layer3_0_aresetn; // @[bfs_remote.scala 229:34]
  wire [31:0] layer3_0_s_axis_tdata; // @[bfs_remote.scala 229:34]
  wire  layer3_0_s_axis_tvalid; // @[bfs_remote.scala 229:34]
  wire [3:0] layer3_0_s_axis_tkeep; // @[bfs_remote.scala 229:34]
  wire  layer3_0_s_axis_tready; // @[bfs_remote.scala 229:34]
  wire  layer3_0_s_axis_tlast; // @[bfs_remote.scala 229:34]
  wire [31:0] layer3_0_m_axis_tdata; // @[bfs_remote.scala 229:34]
  wire  layer3_0_m_axis_tvalid; // @[bfs_remote.scala 229:34]
  wire [3:0] layer3_0_m_axis_tkeep; // @[bfs_remote.scala 229:34]
  wire  layer3_0_m_axis_tready; // @[bfs_remote.scala 229:34]
  wire  layer3_0_m_axis_tlast; // @[bfs_remote.scala 229:34]
  wire  layer3_1_aclk; // @[bfs_remote.scala 229:34]
  wire  layer3_1_aresetn; // @[bfs_remote.scala 229:34]
  wire [31:0] layer3_1_s_axis_tdata; // @[bfs_remote.scala 229:34]
  wire  layer3_1_s_axis_tvalid; // @[bfs_remote.scala 229:34]
  wire [3:0] layer3_1_s_axis_tkeep; // @[bfs_remote.scala 229:34]
  wire  layer3_1_s_axis_tready; // @[bfs_remote.scala 229:34]
  wire  layer3_1_s_axis_tlast; // @[bfs_remote.scala 229:34]
  wire [31:0] layer3_1_m_axis_tdata; // @[bfs_remote.scala 229:34]
  wire  layer3_1_m_axis_tvalid; // @[bfs_remote.scala 229:34]
  wire [3:0] layer3_1_m_axis_tkeep; // @[bfs_remote.scala 229:34]
  wire  layer3_1_m_axis_tready; // @[bfs_remote.scala 229:34]
  wire  layer3_1_m_axis_tlast; // @[bfs_remote.scala 229:34]
  wire  pending_out_aclk; // @[bfs_remote.scala 255:27]
  wire  pending_out_aresetn; // @[bfs_remote.scala 255:27]
  wire [31:0] pending_out_s_axis_tdata; // @[bfs_remote.scala 255:27]
  wire  pending_out_s_axis_tvalid; // @[bfs_remote.scala 255:27]
  wire [3:0] pending_out_s_axis_tkeep; // @[bfs_remote.scala 255:27]
  wire  pending_out_s_axis_tready; // @[bfs_remote.scala 255:27]
  wire  pending_out_s_axis_tlast; // @[bfs_remote.scala 255:27]
  wire [31:0] pending_out_m_axis_tdata; // @[bfs_remote.scala 255:27]
  wire  pending_out_m_axis_tvalid; // @[bfs_remote.scala 255:27]
  wire [3:0] pending_out_m_axis_tkeep; // @[bfs_remote.scala 255:27]
  wire  pending_out_m_axis_tready; // @[bfs_remote.scala 255:27]
  wire  pending_out_m_axis_tlast; // @[bfs_remote.scala 255:27]
  reg [31:0] timing; // @[bfs_remote.scala 184:23]
  wire [31:0] _T_530 = io_period - 32'h3; // @[bfs_remote.scala 186:32]
  wire  _T_531 = timing == _T_530; // @[bfs_remote.scala 186:17]
  wire [31:0] _timing_T_1 = timing + 32'h1; // @[bfs_remote.scala 189:24]
  wire  hittable_0_0 = 4'h0 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE = {{4'd0}, hittable_0_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_0 = 4'h0 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_1 = {{4'd0}, hittable_1_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_1 = _count_WIRE + _count_WIRE_1; // @[bfs_remote.scala 192:97]
  wire  hittable_2_0 = 4'h0 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_2 = {{4'd0}, hittable_2_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_3 = _count_T_1 + _count_WIRE_2; // @[bfs_remote.scala 192:97]
  wire  hittable_3_0 = 4'h0 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_3 = {{4'd0}, hittable_3_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_5 = _count_T_3 + _count_WIRE_3; // @[bfs_remote.scala 192:97]
  wire  hittable_4_0 = 4'h0 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_4 = {{4'd0}, hittable_4_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_7 = _count_T_5 + _count_WIRE_4; // @[bfs_remote.scala 192:97]
  wire  hittable_5_0 = 4'h0 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_5 = {{4'd0}, hittable_5_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_9 = _count_T_7 + _count_WIRE_5; // @[bfs_remote.scala 192:97]
  wire  hittable_6_0 = 4'h0 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_6 = {{4'd0}, hittable_6_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_11 = _count_T_9 + _count_WIRE_6; // @[bfs_remote.scala 192:97]
  wire  hittable_7_0 = 4'h0 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_7 = {{4'd0}, hittable_7_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_13 = _count_T_11 + _count_WIRE_7; // @[bfs_remote.scala 192:97]
  wire  hittable_8_0 = 4'h0 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_8 = {{4'd0}, hittable_8_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_15 = _count_T_13 + _count_WIRE_8; // @[bfs_remote.scala 192:97]
  wire  hittable_9_0 = 4'h0 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_9 = {{4'd0}, hittable_9_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_17 = _count_T_15 + _count_WIRE_9; // @[bfs_remote.scala 192:97]
  wire  hittable_10_0 = 4'h0 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_10 = {{4'd0}, hittable_10_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_19 = _count_T_17 + _count_WIRE_10; // @[bfs_remote.scala 192:97]
  wire  hittable_11_0 = 4'h0 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_11 = {{4'd0}, hittable_11_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_21 = _count_T_19 + _count_WIRE_11; // @[bfs_remote.scala 192:97]
  wire  hittable_12_0 = 4'h0 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_12 = {{4'd0}, hittable_12_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_23 = _count_T_21 + _count_WIRE_12; // @[bfs_remote.scala 192:97]
  wire  hittable_13_0 = 4'h0 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_13 = {{4'd0}, hittable_13_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_25 = _count_T_23 + _count_WIRE_13; // @[bfs_remote.scala 192:97]
  wire  hittable_14_0 = 4'h0 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_14 = {{4'd0}, hittable_14_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_27 = _count_T_25 + _count_WIRE_14; // @[bfs_remote.scala 192:97]
  wire  hittable_15_0 = 4'h0 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_15 = {{4'd0}, hittable_15_0}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_1 = 4'h1 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_16 = {{4'd0}, hittable_0_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_1 = 4'h1 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_17 = {{4'd0}, hittable_1_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_31 = _count_WIRE_16 + _count_WIRE_17; // @[bfs_remote.scala 192:97]
  wire  hittable_2_1 = 4'h1 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_18 = {{4'd0}, hittable_2_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_33 = _count_T_31 + _count_WIRE_18; // @[bfs_remote.scala 192:97]
  wire  hittable_3_1 = 4'h1 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_19 = {{4'd0}, hittable_3_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_35 = _count_T_33 + _count_WIRE_19; // @[bfs_remote.scala 192:97]
  wire  hittable_4_1 = 4'h1 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_20 = {{4'd0}, hittable_4_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_37 = _count_T_35 + _count_WIRE_20; // @[bfs_remote.scala 192:97]
  wire  hittable_5_1 = 4'h1 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_21 = {{4'd0}, hittable_5_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_39 = _count_T_37 + _count_WIRE_21; // @[bfs_remote.scala 192:97]
  wire  hittable_6_1 = 4'h1 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_22 = {{4'd0}, hittable_6_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_41 = _count_T_39 + _count_WIRE_22; // @[bfs_remote.scala 192:97]
  wire  hittable_7_1 = 4'h1 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_23 = {{4'd0}, hittable_7_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_43 = _count_T_41 + _count_WIRE_23; // @[bfs_remote.scala 192:97]
  wire  hittable_8_1 = 4'h1 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_24 = {{4'd0}, hittable_8_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_45 = _count_T_43 + _count_WIRE_24; // @[bfs_remote.scala 192:97]
  wire  hittable_9_1 = 4'h1 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_25 = {{4'd0}, hittable_9_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_47 = _count_T_45 + _count_WIRE_25; // @[bfs_remote.scala 192:97]
  wire  hittable_10_1 = 4'h1 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_26 = {{4'd0}, hittable_10_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_49 = _count_T_47 + _count_WIRE_26; // @[bfs_remote.scala 192:97]
  wire  hittable_11_1 = 4'h1 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_27 = {{4'd0}, hittable_11_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_51 = _count_T_49 + _count_WIRE_27; // @[bfs_remote.scala 192:97]
  wire  hittable_12_1 = 4'h1 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_28 = {{4'd0}, hittable_12_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_53 = _count_T_51 + _count_WIRE_28; // @[bfs_remote.scala 192:97]
  wire  hittable_13_1 = 4'h1 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_29 = {{4'd0}, hittable_13_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_55 = _count_T_53 + _count_WIRE_29; // @[bfs_remote.scala 192:97]
  wire  hittable_14_1 = 4'h1 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_30 = {{4'd0}, hittable_14_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_57 = _count_T_55 + _count_WIRE_30; // @[bfs_remote.scala 192:97]
  wire  hittable_15_1 = 4'h1 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_31 = {{4'd0}, hittable_15_1}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_2 = 4'h2 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_32 = {{4'd0}, hittable_0_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_2 = 4'h2 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_33 = {{4'd0}, hittable_1_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_61 = _count_WIRE_32 + _count_WIRE_33; // @[bfs_remote.scala 192:97]
  wire  hittable_2_2 = 4'h2 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_34 = {{4'd0}, hittable_2_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_63 = _count_T_61 + _count_WIRE_34; // @[bfs_remote.scala 192:97]
  wire  hittable_3_2 = 4'h2 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_35 = {{4'd0}, hittable_3_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_65 = _count_T_63 + _count_WIRE_35; // @[bfs_remote.scala 192:97]
  wire  hittable_4_2 = 4'h2 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_36 = {{4'd0}, hittable_4_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_67 = _count_T_65 + _count_WIRE_36; // @[bfs_remote.scala 192:97]
  wire  hittable_5_2 = 4'h2 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_37 = {{4'd0}, hittable_5_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_69 = _count_T_67 + _count_WIRE_37; // @[bfs_remote.scala 192:97]
  wire  hittable_6_2 = 4'h2 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_38 = {{4'd0}, hittable_6_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_71 = _count_T_69 + _count_WIRE_38; // @[bfs_remote.scala 192:97]
  wire  hittable_7_2 = 4'h2 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_39 = {{4'd0}, hittable_7_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_73 = _count_T_71 + _count_WIRE_39; // @[bfs_remote.scala 192:97]
  wire  hittable_8_2 = 4'h2 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_40 = {{4'd0}, hittable_8_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_75 = _count_T_73 + _count_WIRE_40; // @[bfs_remote.scala 192:97]
  wire  hittable_9_2 = 4'h2 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_41 = {{4'd0}, hittable_9_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_77 = _count_T_75 + _count_WIRE_41; // @[bfs_remote.scala 192:97]
  wire  hittable_10_2 = 4'h2 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_42 = {{4'd0}, hittable_10_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_79 = _count_T_77 + _count_WIRE_42; // @[bfs_remote.scala 192:97]
  wire  hittable_11_2 = 4'h2 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_43 = {{4'd0}, hittable_11_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_81 = _count_T_79 + _count_WIRE_43; // @[bfs_remote.scala 192:97]
  wire  hittable_12_2 = 4'h2 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_44 = {{4'd0}, hittable_12_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_83 = _count_T_81 + _count_WIRE_44; // @[bfs_remote.scala 192:97]
  wire  hittable_13_2 = 4'h2 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_45 = {{4'd0}, hittable_13_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_85 = _count_T_83 + _count_WIRE_45; // @[bfs_remote.scala 192:97]
  wire  hittable_14_2 = 4'h2 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_46 = {{4'd0}, hittable_14_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_87 = _count_T_85 + _count_WIRE_46; // @[bfs_remote.scala 192:97]
  wire  hittable_15_2 = 4'h2 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_47 = {{4'd0}, hittable_15_2}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_3 = 4'h3 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_48 = {{4'd0}, hittable_0_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_3 = 4'h3 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_49 = {{4'd0}, hittable_1_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_91 = _count_WIRE_48 + _count_WIRE_49; // @[bfs_remote.scala 192:97]
  wire  hittable_2_3 = 4'h3 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_50 = {{4'd0}, hittable_2_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_93 = _count_T_91 + _count_WIRE_50; // @[bfs_remote.scala 192:97]
  wire  hittable_3_3 = 4'h3 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_51 = {{4'd0}, hittable_3_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_95 = _count_T_93 + _count_WIRE_51; // @[bfs_remote.scala 192:97]
  wire  hittable_4_3 = 4'h3 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_52 = {{4'd0}, hittable_4_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_97 = _count_T_95 + _count_WIRE_52; // @[bfs_remote.scala 192:97]
  wire  hittable_5_3 = 4'h3 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_53 = {{4'd0}, hittable_5_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_99 = _count_T_97 + _count_WIRE_53; // @[bfs_remote.scala 192:97]
  wire  hittable_6_3 = 4'h3 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_54 = {{4'd0}, hittable_6_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_101 = _count_T_99 + _count_WIRE_54; // @[bfs_remote.scala 192:97]
  wire  hittable_7_3 = 4'h3 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_55 = {{4'd0}, hittable_7_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_103 = _count_T_101 + _count_WIRE_55; // @[bfs_remote.scala 192:97]
  wire  hittable_8_3 = 4'h3 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_56 = {{4'd0}, hittable_8_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_105 = _count_T_103 + _count_WIRE_56; // @[bfs_remote.scala 192:97]
  wire  hittable_9_3 = 4'h3 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_57 = {{4'd0}, hittable_9_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_107 = _count_T_105 + _count_WIRE_57; // @[bfs_remote.scala 192:97]
  wire  hittable_10_3 = 4'h3 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_58 = {{4'd0}, hittable_10_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_109 = _count_T_107 + _count_WIRE_58; // @[bfs_remote.scala 192:97]
  wire  hittable_11_3 = 4'h3 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_59 = {{4'd0}, hittable_11_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_111 = _count_T_109 + _count_WIRE_59; // @[bfs_remote.scala 192:97]
  wire  hittable_12_3 = 4'h3 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_60 = {{4'd0}, hittable_12_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_113 = _count_T_111 + _count_WIRE_60; // @[bfs_remote.scala 192:97]
  wire  hittable_13_3 = 4'h3 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_61 = {{4'd0}, hittable_13_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_115 = _count_T_113 + _count_WIRE_61; // @[bfs_remote.scala 192:97]
  wire  hittable_14_3 = 4'h3 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_62 = {{4'd0}, hittable_14_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_117 = _count_T_115 + _count_WIRE_62; // @[bfs_remote.scala 192:97]
  wire  hittable_15_3 = 4'h3 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_63 = {{4'd0}, hittable_15_3}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_4 = 4'h4 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_64 = {{4'd0}, hittable_0_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_4 = 4'h4 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_65 = {{4'd0}, hittable_1_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_121 = _count_WIRE_64 + _count_WIRE_65; // @[bfs_remote.scala 192:97]
  wire  hittable_2_4 = 4'h4 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_66 = {{4'd0}, hittable_2_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_123 = _count_T_121 + _count_WIRE_66; // @[bfs_remote.scala 192:97]
  wire  hittable_3_4 = 4'h4 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_67 = {{4'd0}, hittable_3_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_125 = _count_T_123 + _count_WIRE_67; // @[bfs_remote.scala 192:97]
  wire  hittable_4_4 = 4'h4 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_68 = {{4'd0}, hittable_4_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_127 = _count_T_125 + _count_WIRE_68; // @[bfs_remote.scala 192:97]
  wire  hittable_5_4 = 4'h4 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_69 = {{4'd0}, hittable_5_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_129 = _count_T_127 + _count_WIRE_69; // @[bfs_remote.scala 192:97]
  wire  hittable_6_4 = 4'h4 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_70 = {{4'd0}, hittable_6_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_131 = _count_T_129 + _count_WIRE_70; // @[bfs_remote.scala 192:97]
  wire  hittable_7_4 = 4'h4 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_71 = {{4'd0}, hittable_7_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_133 = _count_T_131 + _count_WIRE_71; // @[bfs_remote.scala 192:97]
  wire  hittable_8_4 = 4'h4 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_72 = {{4'd0}, hittable_8_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_135 = _count_T_133 + _count_WIRE_72; // @[bfs_remote.scala 192:97]
  wire  hittable_9_4 = 4'h4 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_73 = {{4'd0}, hittable_9_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_137 = _count_T_135 + _count_WIRE_73; // @[bfs_remote.scala 192:97]
  wire  hittable_10_4 = 4'h4 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_74 = {{4'd0}, hittable_10_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_139 = _count_T_137 + _count_WIRE_74; // @[bfs_remote.scala 192:97]
  wire  hittable_11_4 = 4'h4 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_75 = {{4'd0}, hittable_11_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_141 = _count_T_139 + _count_WIRE_75; // @[bfs_remote.scala 192:97]
  wire  hittable_12_4 = 4'h4 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_76 = {{4'd0}, hittable_12_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_143 = _count_T_141 + _count_WIRE_76; // @[bfs_remote.scala 192:97]
  wire  hittable_13_4 = 4'h4 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_77 = {{4'd0}, hittable_13_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_145 = _count_T_143 + _count_WIRE_77; // @[bfs_remote.scala 192:97]
  wire  hittable_14_4 = 4'h4 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_78 = {{4'd0}, hittable_14_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_147 = _count_T_145 + _count_WIRE_78; // @[bfs_remote.scala 192:97]
  wire  hittable_15_4 = 4'h4 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_79 = {{4'd0}, hittable_15_4}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_5 = 4'h5 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_80 = {{4'd0}, hittable_0_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_5 = 4'h5 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_81 = {{4'd0}, hittable_1_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_151 = _count_WIRE_80 + _count_WIRE_81; // @[bfs_remote.scala 192:97]
  wire  hittable_2_5 = 4'h5 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_82 = {{4'd0}, hittable_2_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_153 = _count_T_151 + _count_WIRE_82; // @[bfs_remote.scala 192:97]
  wire  hittable_3_5 = 4'h5 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_83 = {{4'd0}, hittable_3_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_155 = _count_T_153 + _count_WIRE_83; // @[bfs_remote.scala 192:97]
  wire  hittable_4_5 = 4'h5 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_84 = {{4'd0}, hittable_4_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_157 = _count_T_155 + _count_WIRE_84; // @[bfs_remote.scala 192:97]
  wire  hittable_5_5 = 4'h5 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_85 = {{4'd0}, hittable_5_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_159 = _count_T_157 + _count_WIRE_85; // @[bfs_remote.scala 192:97]
  wire  hittable_6_5 = 4'h5 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_86 = {{4'd0}, hittable_6_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_161 = _count_T_159 + _count_WIRE_86; // @[bfs_remote.scala 192:97]
  wire  hittable_7_5 = 4'h5 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_87 = {{4'd0}, hittable_7_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_163 = _count_T_161 + _count_WIRE_87; // @[bfs_remote.scala 192:97]
  wire  hittable_8_5 = 4'h5 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_88 = {{4'd0}, hittable_8_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_165 = _count_T_163 + _count_WIRE_88; // @[bfs_remote.scala 192:97]
  wire  hittable_9_5 = 4'h5 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_89 = {{4'd0}, hittable_9_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_167 = _count_T_165 + _count_WIRE_89; // @[bfs_remote.scala 192:97]
  wire  hittable_10_5 = 4'h5 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_90 = {{4'd0}, hittable_10_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_169 = _count_T_167 + _count_WIRE_90; // @[bfs_remote.scala 192:97]
  wire  hittable_11_5 = 4'h5 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_91 = {{4'd0}, hittable_11_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_171 = _count_T_169 + _count_WIRE_91; // @[bfs_remote.scala 192:97]
  wire  hittable_12_5 = 4'h5 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_92 = {{4'd0}, hittable_12_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_173 = _count_T_171 + _count_WIRE_92; // @[bfs_remote.scala 192:97]
  wire  hittable_13_5 = 4'h5 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_93 = {{4'd0}, hittable_13_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_175 = _count_T_173 + _count_WIRE_93; // @[bfs_remote.scala 192:97]
  wire  hittable_14_5 = 4'h5 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_94 = {{4'd0}, hittable_14_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_177 = _count_T_175 + _count_WIRE_94; // @[bfs_remote.scala 192:97]
  wire  hittable_15_5 = 4'h5 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_95 = {{4'd0}, hittable_15_5}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_6 = 4'h6 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_96 = {{4'd0}, hittable_0_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_6 = 4'h6 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_97 = {{4'd0}, hittable_1_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_181 = _count_WIRE_96 + _count_WIRE_97; // @[bfs_remote.scala 192:97]
  wire  hittable_2_6 = 4'h6 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_98 = {{4'd0}, hittable_2_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_183 = _count_T_181 + _count_WIRE_98; // @[bfs_remote.scala 192:97]
  wire  hittable_3_6 = 4'h6 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_99 = {{4'd0}, hittable_3_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_185 = _count_T_183 + _count_WIRE_99; // @[bfs_remote.scala 192:97]
  wire  hittable_4_6 = 4'h6 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_100 = {{4'd0}, hittable_4_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_187 = _count_T_185 + _count_WIRE_100; // @[bfs_remote.scala 192:97]
  wire  hittable_5_6 = 4'h6 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_101 = {{4'd0}, hittable_5_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_189 = _count_T_187 + _count_WIRE_101; // @[bfs_remote.scala 192:97]
  wire  hittable_6_6 = 4'h6 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_102 = {{4'd0}, hittable_6_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_191 = _count_T_189 + _count_WIRE_102; // @[bfs_remote.scala 192:97]
  wire  hittable_7_6 = 4'h6 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_103 = {{4'd0}, hittable_7_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_193 = _count_T_191 + _count_WIRE_103; // @[bfs_remote.scala 192:97]
  wire  hittable_8_6 = 4'h6 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_104 = {{4'd0}, hittable_8_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_195 = _count_T_193 + _count_WIRE_104; // @[bfs_remote.scala 192:97]
  wire  hittable_9_6 = 4'h6 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_105 = {{4'd0}, hittable_9_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_197 = _count_T_195 + _count_WIRE_105; // @[bfs_remote.scala 192:97]
  wire  hittable_10_6 = 4'h6 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_106 = {{4'd0}, hittable_10_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_199 = _count_T_197 + _count_WIRE_106; // @[bfs_remote.scala 192:97]
  wire  hittable_11_6 = 4'h6 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_107 = {{4'd0}, hittable_11_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_201 = _count_T_199 + _count_WIRE_107; // @[bfs_remote.scala 192:97]
  wire  hittable_12_6 = 4'h6 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_108 = {{4'd0}, hittable_12_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_203 = _count_T_201 + _count_WIRE_108; // @[bfs_remote.scala 192:97]
  wire  hittable_13_6 = 4'h6 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_109 = {{4'd0}, hittable_13_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_205 = _count_T_203 + _count_WIRE_109; // @[bfs_remote.scala 192:97]
  wire  hittable_14_6 = 4'h6 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_110 = {{4'd0}, hittable_14_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_207 = _count_T_205 + _count_WIRE_110; // @[bfs_remote.scala 192:97]
  wire  hittable_15_6 = 4'h6 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_111 = {{4'd0}, hittable_15_6}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_7 = 4'h7 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_112 = {{4'd0}, hittable_0_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_7 = 4'h7 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_113 = {{4'd0}, hittable_1_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_211 = _count_WIRE_112 + _count_WIRE_113; // @[bfs_remote.scala 192:97]
  wire  hittable_2_7 = 4'h7 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_114 = {{4'd0}, hittable_2_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_213 = _count_T_211 + _count_WIRE_114; // @[bfs_remote.scala 192:97]
  wire  hittable_3_7 = 4'h7 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_115 = {{4'd0}, hittable_3_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_215 = _count_T_213 + _count_WIRE_115; // @[bfs_remote.scala 192:97]
  wire  hittable_4_7 = 4'h7 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_116 = {{4'd0}, hittable_4_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_217 = _count_T_215 + _count_WIRE_116; // @[bfs_remote.scala 192:97]
  wire  hittable_5_7 = 4'h7 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_117 = {{4'd0}, hittable_5_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_219 = _count_T_217 + _count_WIRE_117; // @[bfs_remote.scala 192:97]
  wire  hittable_6_7 = 4'h7 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_118 = {{4'd0}, hittable_6_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_221 = _count_T_219 + _count_WIRE_118; // @[bfs_remote.scala 192:97]
  wire  hittable_7_7 = 4'h7 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_119 = {{4'd0}, hittable_7_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_223 = _count_T_221 + _count_WIRE_119; // @[bfs_remote.scala 192:97]
  wire  hittable_8_7 = 4'h7 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_120 = {{4'd0}, hittable_8_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_225 = _count_T_223 + _count_WIRE_120; // @[bfs_remote.scala 192:97]
  wire  hittable_9_7 = 4'h7 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_121 = {{4'd0}, hittable_9_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_227 = _count_T_225 + _count_WIRE_121; // @[bfs_remote.scala 192:97]
  wire  hittable_10_7 = 4'h7 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_122 = {{4'd0}, hittable_10_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_229 = _count_T_227 + _count_WIRE_122; // @[bfs_remote.scala 192:97]
  wire  hittable_11_7 = 4'h7 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_123 = {{4'd0}, hittable_11_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_231 = _count_T_229 + _count_WIRE_123; // @[bfs_remote.scala 192:97]
  wire  hittable_12_7 = 4'h7 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_124 = {{4'd0}, hittable_12_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_233 = _count_T_231 + _count_WIRE_124; // @[bfs_remote.scala 192:97]
  wire  hittable_13_7 = 4'h7 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_125 = {{4'd0}, hittable_13_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_235 = _count_T_233 + _count_WIRE_125; // @[bfs_remote.scala 192:97]
  wire  hittable_14_7 = 4'h7 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_126 = {{4'd0}, hittable_14_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_237 = _count_T_235 + _count_WIRE_126; // @[bfs_remote.scala 192:97]
  wire  hittable_15_7 = 4'h7 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_127 = {{4'd0}, hittable_15_7}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_8 = 4'h8 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_128 = {{4'd0}, hittable_0_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_8 = 4'h8 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_129 = {{4'd0}, hittable_1_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_241 = _count_WIRE_128 + _count_WIRE_129; // @[bfs_remote.scala 192:97]
  wire  hittable_2_8 = 4'h8 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_130 = {{4'd0}, hittable_2_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_243 = _count_T_241 + _count_WIRE_130; // @[bfs_remote.scala 192:97]
  wire  hittable_3_8 = 4'h8 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_131 = {{4'd0}, hittable_3_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_245 = _count_T_243 + _count_WIRE_131; // @[bfs_remote.scala 192:97]
  wire  hittable_4_8 = 4'h8 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_132 = {{4'd0}, hittable_4_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_247 = _count_T_245 + _count_WIRE_132; // @[bfs_remote.scala 192:97]
  wire  hittable_5_8 = 4'h8 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_133 = {{4'd0}, hittable_5_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_249 = _count_T_247 + _count_WIRE_133; // @[bfs_remote.scala 192:97]
  wire  hittable_6_8 = 4'h8 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_134 = {{4'd0}, hittable_6_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_251 = _count_T_249 + _count_WIRE_134; // @[bfs_remote.scala 192:97]
  wire  hittable_7_8 = 4'h8 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_135 = {{4'd0}, hittable_7_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_253 = _count_T_251 + _count_WIRE_135; // @[bfs_remote.scala 192:97]
  wire  hittable_8_8 = 4'h8 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_136 = {{4'd0}, hittable_8_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_255 = _count_T_253 + _count_WIRE_136; // @[bfs_remote.scala 192:97]
  wire  hittable_9_8 = 4'h8 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_137 = {{4'd0}, hittable_9_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_257 = _count_T_255 + _count_WIRE_137; // @[bfs_remote.scala 192:97]
  wire  hittable_10_8 = 4'h8 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_138 = {{4'd0}, hittable_10_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_259 = _count_T_257 + _count_WIRE_138; // @[bfs_remote.scala 192:97]
  wire  hittable_11_8 = 4'h8 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_139 = {{4'd0}, hittable_11_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_261 = _count_T_259 + _count_WIRE_139; // @[bfs_remote.scala 192:97]
  wire  hittable_12_8 = 4'h8 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_140 = {{4'd0}, hittable_12_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_263 = _count_T_261 + _count_WIRE_140; // @[bfs_remote.scala 192:97]
  wire  hittable_13_8 = 4'h8 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_141 = {{4'd0}, hittable_13_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_265 = _count_T_263 + _count_WIRE_141; // @[bfs_remote.scala 192:97]
  wire  hittable_14_8 = 4'h8 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_142 = {{4'd0}, hittable_14_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_267 = _count_T_265 + _count_WIRE_142; // @[bfs_remote.scala 192:97]
  wire  hittable_15_8 = 4'h8 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_143 = {{4'd0}, hittable_15_8}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_9 = 4'h9 == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_144 = {{4'd0}, hittable_0_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_9 = 4'h9 == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_145 = {{4'd0}, hittable_1_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_271 = _count_WIRE_144 + _count_WIRE_145; // @[bfs_remote.scala 192:97]
  wire  hittable_2_9 = 4'h9 == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_146 = {{4'd0}, hittable_2_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_273 = _count_T_271 + _count_WIRE_146; // @[bfs_remote.scala 192:97]
  wire  hittable_3_9 = 4'h9 == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_147 = {{4'd0}, hittable_3_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_275 = _count_T_273 + _count_WIRE_147; // @[bfs_remote.scala 192:97]
  wire  hittable_4_9 = 4'h9 == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_148 = {{4'd0}, hittable_4_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_277 = _count_T_275 + _count_WIRE_148; // @[bfs_remote.scala 192:97]
  wire  hittable_5_9 = 4'h9 == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_149 = {{4'd0}, hittable_5_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_279 = _count_T_277 + _count_WIRE_149; // @[bfs_remote.scala 192:97]
  wire  hittable_6_9 = 4'h9 == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_150 = {{4'd0}, hittable_6_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_281 = _count_T_279 + _count_WIRE_150; // @[bfs_remote.scala 192:97]
  wire  hittable_7_9 = 4'h9 == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_151 = {{4'd0}, hittable_7_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_283 = _count_T_281 + _count_WIRE_151; // @[bfs_remote.scala 192:97]
  wire  hittable_8_9 = 4'h9 == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_152 = {{4'd0}, hittable_8_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_285 = _count_T_283 + _count_WIRE_152; // @[bfs_remote.scala 192:97]
  wire  hittable_9_9 = 4'h9 == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_153 = {{4'd0}, hittable_9_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_287 = _count_T_285 + _count_WIRE_153; // @[bfs_remote.scala 192:97]
  wire  hittable_10_9 = 4'h9 == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_154 = {{4'd0}, hittable_10_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_289 = _count_T_287 + _count_WIRE_154; // @[bfs_remote.scala 192:97]
  wire  hittable_11_9 = 4'h9 == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_155 = {{4'd0}, hittable_11_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_291 = _count_T_289 + _count_WIRE_155; // @[bfs_remote.scala 192:97]
  wire  hittable_12_9 = 4'h9 == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_156 = {{4'd0}, hittable_12_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_293 = _count_T_291 + _count_WIRE_156; // @[bfs_remote.scala 192:97]
  wire  hittable_13_9 = 4'h9 == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_157 = {{4'd0}, hittable_13_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_295 = _count_T_293 + _count_WIRE_157; // @[bfs_remote.scala 192:97]
  wire  hittable_14_9 = 4'h9 == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_158 = {{4'd0}, hittable_14_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_297 = _count_T_295 + _count_WIRE_158; // @[bfs_remote.scala 192:97]
  wire  hittable_15_9 = 4'h9 == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_159 = {{4'd0}, hittable_15_9}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_10 = 4'ha == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_160 = {{4'd0}, hittable_0_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_10 = 4'ha == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_161 = {{4'd0}, hittable_1_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_301 = _count_WIRE_160 + _count_WIRE_161; // @[bfs_remote.scala 192:97]
  wire  hittable_2_10 = 4'ha == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_162 = {{4'd0}, hittable_2_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_303 = _count_T_301 + _count_WIRE_162; // @[bfs_remote.scala 192:97]
  wire  hittable_3_10 = 4'ha == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_163 = {{4'd0}, hittable_3_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_305 = _count_T_303 + _count_WIRE_163; // @[bfs_remote.scala 192:97]
  wire  hittable_4_10 = 4'ha == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_164 = {{4'd0}, hittable_4_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_307 = _count_T_305 + _count_WIRE_164; // @[bfs_remote.scala 192:97]
  wire  hittable_5_10 = 4'ha == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_165 = {{4'd0}, hittable_5_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_309 = _count_T_307 + _count_WIRE_165; // @[bfs_remote.scala 192:97]
  wire  hittable_6_10 = 4'ha == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_166 = {{4'd0}, hittable_6_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_311 = _count_T_309 + _count_WIRE_166; // @[bfs_remote.scala 192:97]
  wire  hittable_7_10 = 4'ha == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_167 = {{4'd0}, hittable_7_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_313 = _count_T_311 + _count_WIRE_167; // @[bfs_remote.scala 192:97]
  wire  hittable_8_10 = 4'ha == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_168 = {{4'd0}, hittable_8_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_315 = _count_T_313 + _count_WIRE_168; // @[bfs_remote.scala 192:97]
  wire  hittable_9_10 = 4'ha == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_169 = {{4'd0}, hittable_9_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_317 = _count_T_315 + _count_WIRE_169; // @[bfs_remote.scala 192:97]
  wire  hittable_10_10 = 4'ha == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_170 = {{4'd0}, hittable_10_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_319 = _count_T_317 + _count_WIRE_170; // @[bfs_remote.scala 192:97]
  wire  hittable_11_10 = 4'ha == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_171 = {{4'd0}, hittable_11_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_321 = _count_T_319 + _count_WIRE_171; // @[bfs_remote.scala 192:97]
  wire  hittable_12_10 = 4'ha == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_172 = {{4'd0}, hittable_12_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_323 = _count_T_321 + _count_WIRE_172; // @[bfs_remote.scala 192:97]
  wire  hittable_13_10 = 4'ha == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_173 = {{4'd0}, hittable_13_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_325 = _count_T_323 + _count_WIRE_173; // @[bfs_remote.scala 192:97]
  wire  hittable_14_10 = 4'ha == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_174 = {{4'd0}, hittable_14_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_327 = _count_T_325 + _count_WIRE_174; // @[bfs_remote.scala 192:97]
  wire  hittable_15_10 = 4'ha == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_175 = {{4'd0}, hittable_15_10}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_11 = 4'hb == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_176 = {{4'd0}, hittable_0_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_11 = 4'hb == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_177 = {{4'd0}, hittable_1_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_331 = _count_WIRE_176 + _count_WIRE_177; // @[bfs_remote.scala 192:97]
  wire  hittable_2_11 = 4'hb == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_178 = {{4'd0}, hittable_2_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_333 = _count_T_331 + _count_WIRE_178; // @[bfs_remote.scala 192:97]
  wire  hittable_3_11 = 4'hb == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_179 = {{4'd0}, hittable_3_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_335 = _count_T_333 + _count_WIRE_179; // @[bfs_remote.scala 192:97]
  wire  hittable_4_11 = 4'hb == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_180 = {{4'd0}, hittable_4_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_337 = _count_T_335 + _count_WIRE_180; // @[bfs_remote.scala 192:97]
  wire  hittable_5_11 = 4'hb == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_181 = {{4'd0}, hittable_5_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_339 = _count_T_337 + _count_WIRE_181; // @[bfs_remote.scala 192:97]
  wire  hittable_6_11 = 4'hb == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_182 = {{4'd0}, hittable_6_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_341 = _count_T_339 + _count_WIRE_182; // @[bfs_remote.scala 192:97]
  wire  hittable_7_11 = 4'hb == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_183 = {{4'd0}, hittable_7_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_343 = _count_T_341 + _count_WIRE_183; // @[bfs_remote.scala 192:97]
  wire  hittable_8_11 = 4'hb == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_184 = {{4'd0}, hittable_8_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_345 = _count_T_343 + _count_WIRE_184; // @[bfs_remote.scala 192:97]
  wire  hittable_9_11 = 4'hb == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_185 = {{4'd0}, hittable_9_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_347 = _count_T_345 + _count_WIRE_185; // @[bfs_remote.scala 192:97]
  wire  hittable_10_11 = 4'hb == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_186 = {{4'd0}, hittable_10_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_349 = _count_T_347 + _count_WIRE_186; // @[bfs_remote.scala 192:97]
  wire  hittable_11_11 = 4'hb == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_187 = {{4'd0}, hittable_11_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_351 = _count_T_349 + _count_WIRE_187; // @[bfs_remote.scala 192:97]
  wire  hittable_12_11 = 4'hb == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_188 = {{4'd0}, hittable_12_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_353 = _count_T_351 + _count_WIRE_188; // @[bfs_remote.scala 192:97]
  wire  hittable_13_11 = 4'hb == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_189 = {{4'd0}, hittable_13_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_355 = _count_T_353 + _count_WIRE_189; // @[bfs_remote.scala 192:97]
  wire  hittable_14_11 = 4'hb == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_190 = {{4'd0}, hittable_14_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_357 = _count_T_355 + _count_WIRE_190; // @[bfs_remote.scala 192:97]
  wire  hittable_15_11 = 4'hb == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_191 = {{4'd0}, hittable_15_11}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_12 = 4'hc == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_192 = {{4'd0}, hittable_0_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_12 = 4'hc == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_193 = {{4'd0}, hittable_1_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_361 = _count_WIRE_192 + _count_WIRE_193; // @[bfs_remote.scala 192:97]
  wire  hittable_2_12 = 4'hc == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_194 = {{4'd0}, hittable_2_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_363 = _count_T_361 + _count_WIRE_194; // @[bfs_remote.scala 192:97]
  wire  hittable_3_12 = 4'hc == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_195 = {{4'd0}, hittable_3_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_365 = _count_T_363 + _count_WIRE_195; // @[bfs_remote.scala 192:97]
  wire  hittable_4_12 = 4'hc == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_196 = {{4'd0}, hittable_4_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_367 = _count_T_365 + _count_WIRE_196; // @[bfs_remote.scala 192:97]
  wire  hittable_5_12 = 4'hc == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_197 = {{4'd0}, hittable_5_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_369 = _count_T_367 + _count_WIRE_197; // @[bfs_remote.scala 192:97]
  wire  hittable_6_12 = 4'hc == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_198 = {{4'd0}, hittable_6_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_371 = _count_T_369 + _count_WIRE_198; // @[bfs_remote.scala 192:97]
  wire  hittable_7_12 = 4'hc == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_199 = {{4'd0}, hittable_7_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_373 = _count_T_371 + _count_WIRE_199; // @[bfs_remote.scala 192:97]
  wire  hittable_8_12 = 4'hc == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_200 = {{4'd0}, hittable_8_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_375 = _count_T_373 + _count_WIRE_200; // @[bfs_remote.scala 192:97]
  wire  hittable_9_12 = 4'hc == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_201 = {{4'd0}, hittable_9_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_377 = _count_T_375 + _count_WIRE_201; // @[bfs_remote.scala 192:97]
  wire  hittable_10_12 = 4'hc == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_202 = {{4'd0}, hittable_10_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_379 = _count_T_377 + _count_WIRE_202; // @[bfs_remote.scala 192:97]
  wire  hittable_11_12 = 4'hc == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_203 = {{4'd0}, hittable_11_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_381 = _count_T_379 + _count_WIRE_203; // @[bfs_remote.scala 192:97]
  wire  hittable_12_12 = 4'hc == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_204 = {{4'd0}, hittable_12_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_383 = _count_T_381 + _count_WIRE_204; // @[bfs_remote.scala 192:97]
  wire  hittable_13_12 = 4'hc == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_205 = {{4'd0}, hittable_13_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_385 = _count_T_383 + _count_WIRE_205; // @[bfs_remote.scala 192:97]
  wire  hittable_14_12 = 4'hc == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_206 = {{4'd0}, hittable_14_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_387 = _count_T_385 + _count_WIRE_206; // @[bfs_remote.scala 192:97]
  wire  hittable_15_12 = 4'hc == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_207 = {{4'd0}, hittable_15_12}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_13 = 4'hd == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_208 = {{4'd0}, hittable_0_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_13 = 4'hd == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_209 = {{4'd0}, hittable_1_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_391 = _count_WIRE_208 + _count_WIRE_209; // @[bfs_remote.scala 192:97]
  wire  hittable_2_13 = 4'hd == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_210 = {{4'd0}, hittable_2_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_393 = _count_T_391 + _count_WIRE_210; // @[bfs_remote.scala 192:97]
  wire  hittable_3_13 = 4'hd == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_211 = {{4'd0}, hittable_3_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_395 = _count_T_393 + _count_WIRE_211; // @[bfs_remote.scala 192:97]
  wire  hittable_4_13 = 4'hd == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_212 = {{4'd0}, hittable_4_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_397 = _count_T_395 + _count_WIRE_212; // @[bfs_remote.scala 192:97]
  wire  hittable_5_13 = 4'hd == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_213 = {{4'd0}, hittable_5_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_399 = _count_T_397 + _count_WIRE_213; // @[bfs_remote.scala 192:97]
  wire  hittable_6_13 = 4'hd == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_214 = {{4'd0}, hittable_6_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_401 = _count_T_399 + _count_WIRE_214; // @[bfs_remote.scala 192:97]
  wire  hittable_7_13 = 4'hd == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_215 = {{4'd0}, hittable_7_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_403 = _count_T_401 + _count_WIRE_215; // @[bfs_remote.scala 192:97]
  wire  hittable_8_13 = 4'hd == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_216 = {{4'd0}, hittable_8_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_405 = _count_T_403 + _count_WIRE_216; // @[bfs_remote.scala 192:97]
  wire  hittable_9_13 = 4'hd == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_217 = {{4'd0}, hittable_9_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_407 = _count_T_405 + _count_WIRE_217; // @[bfs_remote.scala 192:97]
  wire  hittable_10_13 = 4'hd == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_218 = {{4'd0}, hittable_10_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_409 = _count_T_407 + _count_WIRE_218; // @[bfs_remote.scala 192:97]
  wire  hittable_11_13 = 4'hd == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_219 = {{4'd0}, hittable_11_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_411 = _count_T_409 + _count_WIRE_219; // @[bfs_remote.scala 192:97]
  wire  hittable_12_13 = 4'hd == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_220 = {{4'd0}, hittable_12_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_413 = _count_T_411 + _count_WIRE_220; // @[bfs_remote.scala 192:97]
  wire  hittable_13_13 = 4'hd == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_221 = {{4'd0}, hittable_13_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_415 = _count_T_413 + _count_WIRE_221; // @[bfs_remote.scala 192:97]
  wire  hittable_14_13 = 4'hd == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_222 = {{4'd0}, hittable_14_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_417 = _count_T_415 + _count_WIRE_222; // @[bfs_remote.scala 192:97]
  wire  hittable_15_13 = 4'hd == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_223 = {{4'd0}, hittable_15_13}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_14 = 4'he == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_224 = {{4'd0}, hittable_0_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_14 = 4'he == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_225 = {{4'd0}, hittable_1_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_421 = _count_WIRE_224 + _count_WIRE_225; // @[bfs_remote.scala 192:97]
  wire  hittable_2_14 = 4'he == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_226 = {{4'd0}, hittable_2_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_423 = _count_T_421 + _count_WIRE_226; // @[bfs_remote.scala 192:97]
  wire  hittable_3_14 = 4'he == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_227 = {{4'd0}, hittable_3_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_425 = _count_T_423 + _count_WIRE_227; // @[bfs_remote.scala 192:97]
  wire  hittable_4_14 = 4'he == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_228 = {{4'd0}, hittable_4_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_427 = _count_T_425 + _count_WIRE_228; // @[bfs_remote.scala 192:97]
  wire  hittable_5_14 = 4'he == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_229 = {{4'd0}, hittable_5_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_429 = _count_T_427 + _count_WIRE_229; // @[bfs_remote.scala 192:97]
  wire  hittable_6_14 = 4'he == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_230 = {{4'd0}, hittable_6_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_431 = _count_T_429 + _count_WIRE_230; // @[bfs_remote.scala 192:97]
  wire  hittable_7_14 = 4'he == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_231 = {{4'd0}, hittable_7_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_433 = _count_T_431 + _count_WIRE_231; // @[bfs_remote.scala 192:97]
  wire  hittable_8_14 = 4'he == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_232 = {{4'd0}, hittable_8_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_435 = _count_T_433 + _count_WIRE_232; // @[bfs_remote.scala 192:97]
  wire  hittable_9_14 = 4'he == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_233 = {{4'd0}, hittable_9_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_437 = _count_T_435 + _count_WIRE_233; // @[bfs_remote.scala 192:97]
  wire  hittable_10_14 = 4'he == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_234 = {{4'd0}, hittable_10_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_439 = _count_T_437 + _count_WIRE_234; // @[bfs_remote.scala 192:97]
  wire  hittable_11_14 = 4'he == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_235 = {{4'd0}, hittable_11_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_441 = _count_T_439 + _count_WIRE_235; // @[bfs_remote.scala 192:97]
  wire  hittable_12_14 = 4'he == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_236 = {{4'd0}, hittable_12_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_443 = _count_T_441 + _count_WIRE_236; // @[bfs_remote.scala 192:97]
  wire  hittable_13_14 = 4'he == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_237 = {{4'd0}, hittable_13_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_445 = _count_T_443 + _count_WIRE_237; // @[bfs_remote.scala 192:97]
  wire  hittable_14_14 = 4'he == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_238 = {{4'd0}, hittable_14_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_447 = _count_T_445 + _count_WIRE_238; // @[bfs_remote.scala 192:97]
  wire  hittable_15_14 = 4'he == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_239 = {{4'd0}, hittable_15_14}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_0_15 = 4'hf == io_data[5:2] & io_keep[0]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_240 = {{4'd0}, hittable_0_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire  hittable_1_15 = 4'hf == io_data[37:34] & io_keep[1]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_241 = {{4'd0}, hittable_1_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_451 = _count_WIRE_240 + _count_WIRE_241; // @[bfs_remote.scala 192:97]
  wire  hittable_2_15 = 4'hf == io_data[69:66] & io_keep[2]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_242 = {{4'd0}, hittable_2_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_453 = _count_T_451 + _count_WIRE_242; // @[bfs_remote.scala 192:97]
  wire  hittable_3_15 = 4'hf == io_data[101:98] & io_keep[3]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_243 = {{4'd0}, hittable_3_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_455 = _count_T_453 + _count_WIRE_243; // @[bfs_remote.scala 192:97]
  wire  hittable_4_15 = 4'hf == io_data[133:130] & io_keep[4]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_244 = {{4'd0}, hittable_4_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_457 = _count_T_455 + _count_WIRE_244; // @[bfs_remote.scala 192:97]
  wire  hittable_5_15 = 4'hf == io_data[165:162] & io_keep[5]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_245 = {{4'd0}, hittable_5_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_459 = _count_T_457 + _count_WIRE_245; // @[bfs_remote.scala 192:97]
  wire  hittable_6_15 = 4'hf == io_data[197:194] & io_keep[6]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_246 = {{4'd0}, hittable_6_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_461 = _count_T_459 + _count_WIRE_246; // @[bfs_remote.scala 192:97]
  wire  hittable_7_15 = 4'hf == io_data[229:226] & io_keep[7]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_247 = {{4'd0}, hittable_7_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_463 = _count_T_461 + _count_WIRE_247; // @[bfs_remote.scala 192:97]
  wire  hittable_8_15 = 4'hf == io_data[261:258] & io_keep[8]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_248 = {{4'd0}, hittable_8_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_465 = _count_T_463 + _count_WIRE_248; // @[bfs_remote.scala 192:97]
  wire  hittable_9_15 = 4'hf == io_data[293:290] & io_keep[9]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_249 = {{4'd0}, hittable_9_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_467 = _count_T_465 + _count_WIRE_249; // @[bfs_remote.scala 192:97]
  wire  hittable_10_15 = 4'hf == io_data[325:322] & io_keep[10]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_250 = {{4'd0}, hittable_10_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_469 = _count_T_467 + _count_WIRE_250; // @[bfs_remote.scala 192:97]
  wire  hittable_11_15 = 4'hf == io_data[357:354] & io_keep[11]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_251 = {{4'd0}, hittable_11_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_471 = _count_T_469 + _count_WIRE_251; // @[bfs_remote.scala 192:97]
  wire  hittable_12_15 = 4'hf == io_data[389:386] & io_keep[12]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_252 = {{4'd0}, hittable_12_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_473 = _count_T_471 + _count_WIRE_252; // @[bfs_remote.scala 192:97]
  wire  hittable_13_15 = 4'hf == io_data[421:418] & io_keep[13]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_253 = {{4'd0}, hittable_13_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_475 = _count_T_473 + _count_WIRE_253; // @[bfs_remote.scala 192:97]
  wire  hittable_14_15 = 4'hf == io_data[453:450] & io_keep[14]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_254 = {{4'd0}, hittable_14_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  wire [4:0] _count_T_477 = _count_T_475 + _count_WIRE_254; // @[bfs_remote.scala 192:97]
  wire  hittable_15_15 = 4'hf == io_data[485:482] & io_keep[15]; // @[bfs_remote.scala 176:83 bfs_remote.scala 177:26 bfs_remote.scala 179:26]
  wire [4:0] _count_WIRE_255 = {{4'd0}, hittable_15_15}; // @[bfs_remote.scala 192:76 bfs_remote.scala 192:76]
  reg [15:0] count_reg_0; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_1; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_2; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_3; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_4; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_5; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_6; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_7; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_8; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_9; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_10; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_11; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_12; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_13; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_14; // @[bfs_remote.scala 194:26]
  reg [15:0] count_reg_15; // @[bfs_remote.scala 194:26]
  wire [4:0] count_0 = _count_T_27 + _count_WIRE_15; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_294 = {{11'd0}, count_0}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_0_T_1 = count_reg_0 + _GEN_294; // @[bfs_remote.scala 201:20]
  wire [4:0] count_1 = _count_T_57 + _count_WIRE_31; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_295 = {{11'd0}, count_1}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_1_T_1 = count_reg_1 + _GEN_295; // @[bfs_remote.scala 201:20]
  wire [4:0] count_2 = _count_T_87 + _count_WIRE_47; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_296 = {{11'd0}, count_2}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_2_T_1 = count_reg_2 + _GEN_296; // @[bfs_remote.scala 201:20]
  wire [4:0] count_3 = _count_T_117 + _count_WIRE_63; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_297 = {{11'd0}, count_3}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_3_T_1 = count_reg_3 + _GEN_297; // @[bfs_remote.scala 201:20]
  wire [4:0] count_4 = _count_T_147 + _count_WIRE_79; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_298 = {{11'd0}, count_4}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_4_T_1 = count_reg_4 + _GEN_298; // @[bfs_remote.scala 201:20]
  wire [4:0] count_5 = _count_T_177 + _count_WIRE_95; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_299 = {{11'd0}, count_5}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_5_T_1 = count_reg_5 + _GEN_299; // @[bfs_remote.scala 201:20]
  wire [4:0] count_6 = _count_T_207 + _count_WIRE_111; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_300 = {{11'd0}, count_6}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_6_T_1 = count_reg_6 + _GEN_300; // @[bfs_remote.scala 201:20]
  wire [4:0] count_7 = _count_T_237 + _count_WIRE_127; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_301 = {{11'd0}, count_7}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_7_T_1 = count_reg_7 + _GEN_301; // @[bfs_remote.scala 201:20]
  wire [4:0] count_8 = _count_T_267 + _count_WIRE_143; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_302 = {{11'd0}, count_8}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_8_T_1 = count_reg_8 + _GEN_302; // @[bfs_remote.scala 201:20]
  wire [4:0] count_9 = _count_T_297 + _count_WIRE_159; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_303 = {{11'd0}, count_9}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_9_T_1 = count_reg_9 + _GEN_303; // @[bfs_remote.scala 201:20]
  wire [4:0] count_10 = _count_T_327 + _count_WIRE_175; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_304 = {{11'd0}, count_10}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_10_T_1 = count_reg_10 + _GEN_304; // @[bfs_remote.scala 201:20]
  wire [4:0] count_11 = _count_T_357 + _count_WIRE_191; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_305 = {{11'd0}, count_11}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_11_T_1 = count_reg_11 + _GEN_305; // @[bfs_remote.scala 201:20]
  wire [4:0] count_12 = _count_T_387 + _count_WIRE_207; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_306 = {{11'd0}, count_12}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_12_T_1 = count_reg_12 + _GEN_306; // @[bfs_remote.scala 201:20]
  wire [4:0] count_13 = _count_T_417 + _count_WIRE_223; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_307 = {{11'd0}, count_13}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_13_T_1 = count_reg_13 + _GEN_307; // @[bfs_remote.scala 201:20]
  wire [4:0] count_14 = _count_T_447 + _count_WIRE_239; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_308 = {{11'd0}, count_14}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_14_T_1 = count_reg_14 + _GEN_308; // @[bfs_remote.scala 201:20]
  wire [4:0] count_15 = _count_T_477 + _count_WIRE_255; // @[bfs_remote.scala 192:97]
  wire [15:0] _GEN_309 = {{11'd0}, count_15}; // @[bfs_remote.scala 201:20]
  wire [15:0] _count_reg_15_T_1 = count_reg_15 + _GEN_309; // @[bfs_remote.scala 201:20]
  wire [15:0] _layer1_0_io_s_axis_tdata_T_1 = count_reg_0 > count_reg_1 ? count_reg_0 : count_reg_1; // @[bfs_remote.scala 213:31]
  wire [15:0] _layer1_1_io_s_axis_tdata_T_1 = count_reg_2 > count_reg_3 ? count_reg_2 : count_reg_3; // @[bfs_remote.scala 213:31]
  wire [15:0] _layer1_2_io_s_axis_tdata_T_1 = count_reg_4 > count_reg_5 ? count_reg_4 : count_reg_5; // @[bfs_remote.scala 213:31]
  wire [15:0] _layer1_3_io_s_axis_tdata_T_1 = count_reg_6 > count_reg_7 ? count_reg_6 : count_reg_7; // @[bfs_remote.scala 213:31]
  wire [15:0] _layer1_4_io_s_axis_tdata_T_1 = count_reg_8 > count_reg_9 ? count_reg_8 : count_reg_9; // @[bfs_remote.scala 213:31]
  wire [15:0] _layer1_5_io_s_axis_tdata_T_1 = count_reg_10 > count_reg_11 ? count_reg_10 : count_reg_11; // @[bfs_remote.scala 213:31]
  wire [15:0] _layer1_6_io_s_axis_tdata_T_1 = count_reg_12 > count_reg_13 ? count_reg_12 : count_reg_13; // @[bfs_remote.scala 213:31]
  wire [15:0] _layer1_7_io_s_axis_tdata_T_1 = count_reg_14 > count_reg_15 ? count_reg_14 : count_reg_15; // @[bfs_remote.scala 213:31]
  wire [31:0] max_a = layer3_0_m_axis_tdata > layer3_1_m_axis_tdata ? layer3_0_m_axis_tdata : layer3_1_m_axis_tdata; // @[bfs_remote.scala 241:18]
  wire [16:0] _GEN_310 = {max_a[15:0], 1'h0}; // @[bfs_remote.scala 251:37]
  wire [30:0] pending_options_1 = {{14'd0}, _GEN_310}; // @[bfs_remote.scala 251:37]
  wire [30:0] _GEN_312 = {{11'd0}, max_a[19:0]}; // @[bfs_remote.scala 249:69]
  wire [30:0] pending_options_2 = pending_options_1 + _GEN_312; // @[bfs_remote.scala 249:69]
  wire [17:0] _GEN_313 = {max_a[15:0], 2'h0}; // @[bfs_remote.scala 251:37]
  wire [30:0] pending_options_3 = {{13'd0}, _GEN_313}; // @[bfs_remote.scala 251:37]
  wire [2:0] _GEN_314 = {{1'd0}, io_idol_fpga_num}; // @[bfs_remote.scala 258:61]
  wire [2:0] _pending_out_io_s_axis_tdata_T_1 = 3'h4 - _GEN_314; // @[bfs_remote.scala 258:61]
  wire [2:0] _pending_out_io_s_axis_tdata_T_3 = _pending_out_io_s_axis_tdata_T_1 - 3'h1; // @[bfs_remote.scala 258:80]
  wire [30:0] _GEN_291 = 2'h1 == _pending_out_io_s_axis_tdata_T_3[1:0] ? pending_options_1 : _GEN_312; // @[bfs_remote.scala 258:87 bfs_remote.scala 258:87]
  wire [30:0] _GEN_292 = 2'h2 == _pending_out_io_s_axis_tdata_T_3[1:0] ? pending_options_2 : _GEN_291; // @[bfs_remote.scala 258:87 bfs_remote.scala 258:87]
  wire [30:0] _GEN_293 = 2'h3 == _pending_out_io_s_axis_tdata_T_3[1:0] ? pending_options_3 : _GEN_292; // @[bfs_remote.scala 258:87 bfs_remote.scala 258:87]
  wire [31:0] _GEN_315 = {{1'd0}, _GEN_293}; // @[bfs_remote.scala 258:87]
  flow_control_reg layer1_0 ( // @[bfs_remote.scala 208:34]
    .aclk(layer1_0_aclk),
    .aresetn(layer1_0_aresetn),
    .s_axis_tdata(layer1_0_s_axis_tdata),
    .s_axis_tvalid(layer1_0_s_axis_tvalid),
    .s_axis_tkeep(layer1_0_s_axis_tkeep),
    .s_axis_tready(layer1_0_s_axis_tready),
    .s_axis_tlast(layer1_0_s_axis_tlast),
    .m_axis_tdata(layer1_0_m_axis_tdata),
    .m_axis_tvalid(layer1_0_m_axis_tvalid),
    .m_axis_tkeep(layer1_0_m_axis_tkeep),
    .m_axis_tready(layer1_0_m_axis_tready),
    .m_axis_tlast(layer1_0_m_axis_tlast)
  );
  flow_control_reg layer1_1 ( // @[bfs_remote.scala 208:34]
    .aclk(layer1_1_aclk),
    .aresetn(layer1_1_aresetn),
    .s_axis_tdata(layer1_1_s_axis_tdata),
    .s_axis_tvalid(layer1_1_s_axis_tvalid),
    .s_axis_tkeep(layer1_1_s_axis_tkeep),
    .s_axis_tready(layer1_1_s_axis_tready),
    .s_axis_tlast(layer1_1_s_axis_tlast),
    .m_axis_tdata(layer1_1_m_axis_tdata),
    .m_axis_tvalid(layer1_1_m_axis_tvalid),
    .m_axis_tkeep(layer1_1_m_axis_tkeep),
    .m_axis_tready(layer1_1_m_axis_tready),
    .m_axis_tlast(layer1_1_m_axis_tlast)
  );
  flow_control_reg layer1_2 ( // @[bfs_remote.scala 208:34]
    .aclk(layer1_2_aclk),
    .aresetn(layer1_2_aresetn),
    .s_axis_tdata(layer1_2_s_axis_tdata),
    .s_axis_tvalid(layer1_2_s_axis_tvalid),
    .s_axis_tkeep(layer1_2_s_axis_tkeep),
    .s_axis_tready(layer1_2_s_axis_tready),
    .s_axis_tlast(layer1_2_s_axis_tlast),
    .m_axis_tdata(layer1_2_m_axis_tdata),
    .m_axis_tvalid(layer1_2_m_axis_tvalid),
    .m_axis_tkeep(layer1_2_m_axis_tkeep),
    .m_axis_tready(layer1_2_m_axis_tready),
    .m_axis_tlast(layer1_2_m_axis_tlast)
  );
  flow_control_reg layer1_3 ( // @[bfs_remote.scala 208:34]
    .aclk(layer1_3_aclk),
    .aresetn(layer1_3_aresetn),
    .s_axis_tdata(layer1_3_s_axis_tdata),
    .s_axis_tvalid(layer1_3_s_axis_tvalid),
    .s_axis_tkeep(layer1_3_s_axis_tkeep),
    .s_axis_tready(layer1_3_s_axis_tready),
    .s_axis_tlast(layer1_3_s_axis_tlast),
    .m_axis_tdata(layer1_3_m_axis_tdata),
    .m_axis_tvalid(layer1_3_m_axis_tvalid),
    .m_axis_tkeep(layer1_3_m_axis_tkeep),
    .m_axis_tready(layer1_3_m_axis_tready),
    .m_axis_tlast(layer1_3_m_axis_tlast)
  );
  flow_control_reg layer1_4 ( // @[bfs_remote.scala 208:34]
    .aclk(layer1_4_aclk),
    .aresetn(layer1_4_aresetn),
    .s_axis_tdata(layer1_4_s_axis_tdata),
    .s_axis_tvalid(layer1_4_s_axis_tvalid),
    .s_axis_tkeep(layer1_4_s_axis_tkeep),
    .s_axis_tready(layer1_4_s_axis_tready),
    .s_axis_tlast(layer1_4_s_axis_tlast),
    .m_axis_tdata(layer1_4_m_axis_tdata),
    .m_axis_tvalid(layer1_4_m_axis_tvalid),
    .m_axis_tkeep(layer1_4_m_axis_tkeep),
    .m_axis_tready(layer1_4_m_axis_tready),
    .m_axis_tlast(layer1_4_m_axis_tlast)
  );
  flow_control_reg layer1_5 ( // @[bfs_remote.scala 208:34]
    .aclk(layer1_5_aclk),
    .aresetn(layer1_5_aresetn),
    .s_axis_tdata(layer1_5_s_axis_tdata),
    .s_axis_tvalid(layer1_5_s_axis_tvalid),
    .s_axis_tkeep(layer1_5_s_axis_tkeep),
    .s_axis_tready(layer1_5_s_axis_tready),
    .s_axis_tlast(layer1_5_s_axis_tlast),
    .m_axis_tdata(layer1_5_m_axis_tdata),
    .m_axis_tvalid(layer1_5_m_axis_tvalid),
    .m_axis_tkeep(layer1_5_m_axis_tkeep),
    .m_axis_tready(layer1_5_m_axis_tready),
    .m_axis_tlast(layer1_5_m_axis_tlast)
  );
  flow_control_reg layer1_6 ( // @[bfs_remote.scala 208:34]
    .aclk(layer1_6_aclk),
    .aresetn(layer1_6_aresetn),
    .s_axis_tdata(layer1_6_s_axis_tdata),
    .s_axis_tvalid(layer1_6_s_axis_tvalid),
    .s_axis_tkeep(layer1_6_s_axis_tkeep),
    .s_axis_tready(layer1_6_s_axis_tready),
    .s_axis_tlast(layer1_6_s_axis_tlast),
    .m_axis_tdata(layer1_6_m_axis_tdata),
    .m_axis_tvalid(layer1_6_m_axis_tvalid),
    .m_axis_tkeep(layer1_6_m_axis_tkeep),
    .m_axis_tready(layer1_6_m_axis_tready),
    .m_axis_tlast(layer1_6_m_axis_tlast)
  );
  flow_control_reg layer1_7 ( // @[bfs_remote.scala 208:34]
    .aclk(layer1_7_aclk),
    .aresetn(layer1_7_aresetn),
    .s_axis_tdata(layer1_7_s_axis_tdata),
    .s_axis_tvalid(layer1_7_s_axis_tvalid),
    .s_axis_tkeep(layer1_7_s_axis_tkeep),
    .s_axis_tready(layer1_7_s_axis_tready),
    .s_axis_tlast(layer1_7_s_axis_tlast),
    .m_axis_tdata(layer1_7_m_axis_tdata),
    .m_axis_tvalid(layer1_7_m_axis_tvalid),
    .m_axis_tkeep(layer1_7_m_axis_tkeep),
    .m_axis_tready(layer1_7_m_axis_tready),
    .m_axis_tlast(layer1_7_m_axis_tlast)
  );
  flow_control_reg layer2_0 ( // @[bfs_remote.scala 217:34]
    .aclk(layer2_0_aclk),
    .aresetn(layer2_0_aresetn),
    .s_axis_tdata(layer2_0_s_axis_tdata),
    .s_axis_tvalid(layer2_0_s_axis_tvalid),
    .s_axis_tkeep(layer2_0_s_axis_tkeep),
    .s_axis_tready(layer2_0_s_axis_tready),
    .s_axis_tlast(layer2_0_s_axis_tlast),
    .m_axis_tdata(layer2_0_m_axis_tdata),
    .m_axis_tvalid(layer2_0_m_axis_tvalid),
    .m_axis_tkeep(layer2_0_m_axis_tkeep),
    .m_axis_tready(layer2_0_m_axis_tready),
    .m_axis_tlast(layer2_0_m_axis_tlast)
  );
  flow_control_reg layer2_1 ( // @[bfs_remote.scala 217:34]
    .aclk(layer2_1_aclk),
    .aresetn(layer2_1_aresetn),
    .s_axis_tdata(layer2_1_s_axis_tdata),
    .s_axis_tvalid(layer2_1_s_axis_tvalid),
    .s_axis_tkeep(layer2_1_s_axis_tkeep),
    .s_axis_tready(layer2_1_s_axis_tready),
    .s_axis_tlast(layer2_1_s_axis_tlast),
    .m_axis_tdata(layer2_1_m_axis_tdata),
    .m_axis_tvalid(layer2_1_m_axis_tvalid),
    .m_axis_tkeep(layer2_1_m_axis_tkeep),
    .m_axis_tready(layer2_1_m_axis_tready),
    .m_axis_tlast(layer2_1_m_axis_tlast)
  );
  flow_control_reg layer2_2 ( // @[bfs_remote.scala 217:34]
    .aclk(layer2_2_aclk),
    .aresetn(layer2_2_aresetn),
    .s_axis_tdata(layer2_2_s_axis_tdata),
    .s_axis_tvalid(layer2_2_s_axis_tvalid),
    .s_axis_tkeep(layer2_2_s_axis_tkeep),
    .s_axis_tready(layer2_2_s_axis_tready),
    .s_axis_tlast(layer2_2_s_axis_tlast),
    .m_axis_tdata(layer2_2_m_axis_tdata),
    .m_axis_tvalid(layer2_2_m_axis_tvalid),
    .m_axis_tkeep(layer2_2_m_axis_tkeep),
    .m_axis_tready(layer2_2_m_axis_tready),
    .m_axis_tlast(layer2_2_m_axis_tlast)
  );
  flow_control_reg layer2_3 ( // @[bfs_remote.scala 217:34]
    .aclk(layer2_3_aclk),
    .aresetn(layer2_3_aresetn),
    .s_axis_tdata(layer2_3_s_axis_tdata),
    .s_axis_tvalid(layer2_3_s_axis_tvalid),
    .s_axis_tkeep(layer2_3_s_axis_tkeep),
    .s_axis_tready(layer2_3_s_axis_tready),
    .s_axis_tlast(layer2_3_s_axis_tlast),
    .m_axis_tdata(layer2_3_m_axis_tdata),
    .m_axis_tvalid(layer2_3_m_axis_tvalid),
    .m_axis_tkeep(layer2_3_m_axis_tkeep),
    .m_axis_tready(layer2_3_m_axis_tready),
    .m_axis_tlast(layer2_3_m_axis_tlast)
  );
  flow_control_reg layer3_0 ( // @[bfs_remote.scala 229:34]
    .aclk(layer3_0_aclk),
    .aresetn(layer3_0_aresetn),
    .s_axis_tdata(layer3_0_s_axis_tdata),
    .s_axis_tvalid(layer3_0_s_axis_tvalid),
    .s_axis_tkeep(layer3_0_s_axis_tkeep),
    .s_axis_tready(layer3_0_s_axis_tready),
    .s_axis_tlast(layer3_0_s_axis_tlast),
    .m_axis_tdata(layer3_0_m_axis_tdata),
    .m_axis_tvalid(layer3_0_m_axis_tvalid),
    .m_axis_tkeep(layer3_0_m_axis_tkeep),
    .m_axis_tready(layer3_0_m_axis_tready),
    .m_axis_tlast(layer3_0_m_axis_tlast)
  );
  flow_control_reg layer3_1 ( // @[bfs_remote.scala 229:34]
    .aclk(layer3_1_aclk),
    .aresetn(layer3_1_aresetn),
    .s_axis_tdata(layer3_1_s_axis_tdata),
    .s_axis_tvalid(layer3_1_s_axis_tvalid),
    .s_axis_tkeep(layer3_1_s_axis_tkeep),
    .s_axis_tready(layer3_1_s_axis_tready),
    .s_axis_tlast(layer3_1_s_axis_tlast),
    .m_axis_tdata(layer3_1_m_axis_tdata),
    .m_axis_tvalid(layer3_1_m_axis_tvalid),
    .m_axis_tkeep(layer3_1_m_axis_tkeep),
    .m_axis_tready(layer3_1_m_axis_tready),
    .m_axis_tlast(layer3_1_m_axis_tlast)
  );
  flow_control_reg pending_out ( // @[bfs_remote.scala 255:27]
    .aclk(pending_out_aclk),
    .aresetn(pending_out_aresetn),
    .s_axis_tdata(pending_out_s_axis_tdata),
    .s_axis_tvalid(pending_out_s_axis_tvalid),
    .s_axis_tkeep(pending_out_s_axis_tkeep),
    .s_axis_tready(pending_out_s_axis_tready),
    .s_axis_tlast(pending_out_s_axis_tlast),
    .m_axis_tdata(pending_out_m_axis_tdata),
    .m_axis_tvalid(pending_out_m_axis_tvalid),
    .m_axis_tkeep(pending_out_m_axis_tkeep),
    .m_axis_tready(pending_out_m_axis_tready),
    .m_axis_tlast(pending_out_m_axis_tlast)
  );
  assign io_pending_valid = pending_out_m_axis_tvalid & pending_out_m_axis_tready; // @[bfs_remote.scala 264:52]
  assign io_pending_bits = pending_out_m_axis_tdata; // @[bfs_remote.scala 263:19]
  assign layer1_0_aclk = clock; // @[bfs_remote.scala 211:32]
  assign layer1_0_aresetn = ~reset; // @[bfs_remote.scala 212:23]
  assign layer1_0_s_axis_tdata = {{16'd0}, _layer1_0_io_s_axis_tdata_T_1}; // @[bfs_remote.scala 213:31]
  assign layer1_0_s_axis_tvalid = _T_531 & io_handshake & io_handshake_last; // @[bfs_remote.scala 214:74]
  assign layer1_0_s_axis_tkeep = 4'h0;
  assign layer1_0_s_axis_tlast = 1'h0;
  assign layer1_0_m_axis_tready = layer2_0_s_axis_tready; // @[bfs_remote.scala 225:36]
  assign layer1_1_aclk = clock; // @[bfs_remote.scala 211:32]
  assign layer1_1_aresetn = ~reset; // @[bfs_remote.scala 212:23]
  assign layer1_1_s_axis_tdata = {{16'd0}, _layer1_1_io_s_axis_tdata_T_1}; // @[bfs_remote.scala 213:31]
  assign layer1_1_s_axis_tvalid = _T_531 & io_handshake & io_handshake_last; // @[bfs_remote.scala 214:74]
  assign layer1_1_s_axis_tkeep = 4'h0;
  assign layer1_1_s_axis_tlast = 1'h0;
  assign layer1_1_m_axis_tready = layer2_0_s_axis_tready; // @[bfs_remote.scala 226:38]
  assign layer1_2_aclk = clock; // @[bfs_remote.scala 211:32]
  assign layer1_2_aresetn = ~reset; // @[bfs_remote.scala 212:23]
  assign layer1_2_s_axis_tdata = {{16'd0}, _layer1_2_io_s_axis_tdata_T_1}; // @[bfs_remote.scala 213:31]
  assign layer1_2_s_axis_tvalid = _T_531 & io_handshake & io_handshake_last; // @[bfs_remote.scala 214:74]
  assign layer1_2_s_axis_tkeep = 4'h0;
  assign layer1_2_s_axis_tlast = 1'h0;
  assign layer1_2_m_axis_tready = layer2_1_s_axis_tready; // @[bfs_remote.scala 225:36]
  assign layer1_3_aclk = clock; // @[bfs_remote.scala 211:32]
  assign layer1_3_aresetn = ~reset; // @[bfs_remote.scala 212:23]
  assign layer1_3_s_axis_tdata = {{16'd0}, _layer1_3_io_s_axis_tdata_T_1}; // @[bfs_remote.scala 213:31]
  assign layer1_3_s_axis_tvalid = _T_531 & io_handshake & io_handshake_last; // @[bfs_remote.scala 214:74]
  assign layer1_3_s_axis_tkeep = 4'h0;
  assign layer1_3_s_axis_tlast = 1'h0;
  assign layer1_3_m_axis_tready = layer2_1_s_axis_tready; // @[bfs_remote.scala 226:38]
  assign layer1_4_aclk = clock; // @[bfs_remote.scala 211:32]
  assign layer1_4_aresetn = ~reset; // @[bfs_remote.scala 212:23]
  assign layer1_4_s_axis_tdata = {{16'd0}, _layer1_4_io_s_axis_tdata_T_1}; // @[bfs_remote.scala 213:31]
  assign layer1_4_s_axis_tvalid = _T_531 & io_handshake & io_handshake_last; // @[bfs_remote.scala 214:74]
  assign layer1_4_s_axis_tkeep = 4'h0;
  assign layer1_4_s_axis_tlast = 1'h0;
  assign layer1_4_m_axis_tready = layer2_2_s_axis_tready; // @[bfs_remote.scala 225:36]
  assign layer1_5_aclk = clock; // @[bfs_remote.scala 211:32]
  assign layer1_5_aresetn = ~reset; // @[bfs_remote.scala 212:23]
  assign layer1_5_s_axis_tdata = {{16'd0}, _layer1_5_io_s_axis_tdata_T_1}; // @[bfs_remote.scala 213:31]
  assign layer1_5_s_axis_tvalid = _T_531 & io_handshake & io_handshake_last; // @[bfs_remote.scala 214:74]
  assign layer1_5_s_axis_tkeep = 4'h0;
  assign layer1_5_s_axis_tlast = 1'h0;
  assign layer1_5_m_axis_tready = layer2_2_s_axis_tready; // @[bfs_remote.scala 226:38]
  assign layer1_6_aclk = clock; // @[bfs_remote.scala 211:32]
  assign layer1_6_aresetn = ~reset; // @[bfs_remote.scala 212:23]
  assign layer1_6_s_axis_tdata = {{16'd0}, _layer1_6_io_s_axis_tdata_T_1}; // @[bfs_remote.scala 213:31]
  assign layer1_6_s_axis_tvalid = _T_531 & io_handshake & io_handshake_last; // @[bfs_remote.scala 214:74]
  assign layer1_6_s_axis_tkeep = 4'h0;
  assign layer1_6_s_axis_tlast = 1'h0;
  assign layer1_6_m_axis_tready = layer2_3_s_axis_tready; // @[bfs_remote.scala 225:36]
  assign layer1_7_aclk = clock; // @[bfs_remote.scala 211:32]
  assign layer1_7_aresetn = ~reset; // @[bfs_remote.scala 212:23]
  assign layer1_7_s_axis_tdata = {{16'd0}, _layer1_7_io_s_axis_tdata_T_1}; // @[bfs_remote.scala 213:31]
  assign layer1_7_s_axis_tvalid = _T_531 & io_handshake & io_handshake_last; // @[bfs_remote.scala 214:74]
  assign layer1_7_s_axis_tkeep = 4'h0;
  assign layer1_7_s_axis_tlast = 1'h0;
  assign layer1_7_m_axis_tready = layer2_3_s_axis_tready; // @[bfs_remote.scala 226:38]
  assign layer2_0_aclk = clock; // @[bfs_remote.scala 220:32]
  assign layer2_0_aresetn = ~reset; // @[bfs_remote.scala 221:23]
  assign layer2_0_s_axis_tdata = layer1_0_m_axis_tdata > layer1_1_m_axis_tdata ? layer1_0_m_axis_tdata :
    layer1_1_m_axis_tdata; // @[bfs_remote.scala 222:31]
  assign layer2_0_s_axis_tvalid = layer1_0_m_axis_tvalid & layer1_1_m_axis_tvalid; // @[bfs_remote.scala 224:58]
  assign layer2_0_s_axis_tkeep = 4'h0;
  assign layer2_0_s_axis_tlast = 1'h0;
  assign layer2_0_m_axis_tready = layer3_0_s_axis_tready; // @[bfs_remote.scala 237:36]
  assign layer2_1_aclk = clock; // @[bfs_remote.scala 220:32]
  assign layer2_1_aresetn = ~reset; // @[bfs_remote.scala 221:23]
  assign layer2_1_s_axis_tdata = layer1_2_m_axis_tdata > layer1_3_m_axis_tdata ? layer1_2_m_axis_tdata :
    layer1_3_m_axis_tdata; // @[bfs_remote.scala 222:31]
  assign layer2_1_s_axis_tvalid = layer1_2_m_axis_tvalid & layer1_3_m_axis_tvalid; // @[bfs_remote.scala 224:58]
  assign layer2_1_s_axis_tkeep = 4'h0;
  assign layer2_1_s_axis_tlast = 1'h0;
  assign layer2_1_m_axis_tready = layer3_0_s_axis_tready; // @[bfs_remote.scala 238:38]
  assign layer2_2_aclk = clock; // @[bfs_remote.scala 220:32]
  assign layer2_2_aresetn = ~reset; // @[bfs_remote.scala 221:23]
  assign layer2_2_s_axis_tdata = layer1_4_m_axis_tdata > layer1_5_m_axis_tdata ? layer1_4_m_axis_tdata :
    layer1_5_m_axis_tdata; // @[bfs_remote.scala 222:31]
  assign layer2_2_s_axis_tvalid = layer1_4_m_axis_tvalid & layer1_5_m_axis_tvalid; // @[bfs_remote.scala 224:58]
  assign layer2_2_s_axis_tkeep = 4'h0;
  assign layer2_2_s_axis_tlast = 1'h0;
  assign layer2_2_m_axis_tready = layer3_1_s_axis_tready; // @[bfs_remote.scala 237:36]
  assign layer2_3_aclk = clock; // @[bfs_remote.scala 220:32]
  assign layer2_3_aresetn = ~reset; // @[bfs_remote.scala 221:23]
  assign layer2_3_s_axis_tdata = layer1_6_m_axis_tdata > layer1_7_m_axis_tdata ? layer1_6_m_axis_tdata :
    layer1_7_m_axis_tdata; // @[bfs_remote.scala 222:31]
  assign layer2_3_s_axis_tvalid = layer1_6_m_axis_tvalid & layer1_7_m_axis_tvalid; // @[bfs_remote.scala 224:58]
  assign layer2_3_s_axis_tkeep = 4'h0;
  assign layer2_3_s_axis_tlast = 1'h0;
  assign layer2_3_m_axis_tready = layer3_1_s_axis_tready; // @[bfs_remote.scala 238:38]
  assign layer3_0_aclk = clock; // @[bfs_remote.scala 232:32]
  assign layer3_0_aresetn = ~reset; // @[bfs_remote.scala 233:23]
  assign layer3_0_s_axis_tdata = layer2_0_m_axis_tdata > layer2_1_m_axis_tdata ? layer2_0_m_axis_tdata :
    layer2_1_m_axis_tdata; // @[bfs_remote.scala 234:31]
  assign layer3_0_s_axis_tvalid = layer2_0_m_axis_tvalid & layer2_1_m_axis_tvalid; // @[bfs_remote.scala 236:58]
  assign layer3_0_s_axis_tkeep = 4'h0;
  assign layer3_0_s_axis_tlast = 1'h0;
  assign layer3_0_m_axis_tready = pending_out_s_axis_tready; // @[bfs_remote.scala 260:30]
  assign layer3_1_aclk = clock; // @[bfs_remote.scala 232:32]
  assign layer3_1_aresetn = ~reset; // @[bfs_remote.scala 233:23]
  assign layer3_1_s_axis_tdata = layer2_2_m_axis_tdata > layer2_3_m_axis_tdata ? layer2_2_m_axis_tdata :
    layer2_3_m_axis_tdata; // @[bfs_remote.scala 234:31]
  assign layer3_1_s_axis_tvalid = layer2_2_m_axis_tvalid & layer2_3_m_axis_tvalid; // @[bfs_remote.scala 236:58]
  assign layer3_1_s_axis_tkeep = 4'h0;
  assign layer3_1_s_axis_tlast = 1'h0;
  assign layer3_1_m_axis_tready = pending_out_s_axis_tready; // @[bfs_remote.scala 261:30]
  assign pending_out_aclk = clock; // @[bfs_remote.scala 256:38]
  assign pending_out_aresetn = ~reset; // @[bfs_remote.scala 257:29]
  assign pending_out_s_axis_tdata = _GEN_315 - io_parameter; // @[bfs_remote.scala 258:87]
  assign pending_out_s_axis_tvalid = layer3_0_m_axis_tvalid & layer3_1_m_axis_tvalid; // @[bfs_remote.scala 259:62]
  assign pending_out_s_axis_tkeep = 4'h0;
  assign pending_out_s_axis_tlast = 1'h0;
  assign pending_out_m_axis_tready = io_handshake & io_handshake_last; // @[bfs_remote.scala 265:48]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 184:23]
      timing <= 32'h0; // @[bfs_remote.scala 184:23]
    end else if (io_handshake & io_handshake_last) begin // @[bfs_remote.scala 185:42]
      if (timing == _T_530) begin // @[bfs_remote.scala 186:39]
        timing <= 32'h0; // @[bfs_remote.scala 187:14]
      end else begin
        timing <= _timing_T_1; // @[bfs_remote.scala 189:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_0 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_0 <= {{11'd0}, count_0}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_0 <= _count_reg_0_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_1 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_1 <= {{11'd0}, count_1}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_1 <= _count_reg_1_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_2 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_2 <= {{11'd0}, count_2}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_2 <= _count_reg_2_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_3 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_3 <= {{11'd0}, count_3}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_3 <= _count_reg_3_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_4 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_4 <= {{11'd0}, count_4}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_4 <= _count_reg_4_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_5 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_5 <= {{11'd0}, count_5}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_5 <= _count_reg_5_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_6 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_6 <= {{11'd0}, count_6}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_6 <= _count_reg_6_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_7 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_7 <= {{11'd0}, count_7}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_7 <= _count_reg_7_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_8 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_8 <= {{11'd0}, count_8}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_8 <= _count_reg_8_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_9 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_9 <= {{11'd0}, count_9}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_9 <= _count_reg_9_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_10 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_10 <= {{11'd0}, count_10}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_10 <= _count_reg_10_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_11 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_11 <= {{11'd0}, count_11}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_11 <= _count_reg_11_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_12 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_12 <= {{11'd0}, count_12}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_12 <= _count_reg_12_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_13 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_13 <= {{11'd0}, count_13}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_13 <= _count_reg_13_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_14 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_14 <= {{11'd0}, count_14}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_14 <= _count_reg_14_T_1; // @[bfs_remote.scala 201:14]
      end
    end
    if (reset) begin // @[bfs_remote.scala 194:26]
      count_reg_15 <= 16'h0; // @[bfs_remote.scala 194:26]
    end else if (io_handshake) begin // @[bfs_remote.scala 197:25]
      if (_T_531 & io_handshake_last) begin // @[bfs_remote.scala 198:64]
        count_reg_15 <= {{11'd0}, count_15}; // @[bfs_remote.scala 199:14]
      end else begin
        count_reg_15 <= _count_reg_15_T_1; // @[bfs_remote.scala 201:14]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  timing = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  count_reg_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  count_reg_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  count_reg_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  count_reg_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  count_reg_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  count_reg_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  count_reg_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  count_reg_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  count_reg_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  count_reg_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  count_reg_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  count_reg_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  count_reg_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  count_reg_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  count_reg_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  count_reg_15 = _RAND_16[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Remote_Apply(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_remote_out_ready,
  output         io_remote_out_valid,
  output [511:0] io_remote_out_bits_tdata,
  output [63:0]  io_remote_out_bits_tkeep,
  output         io_remote_out_bits_tlast,
  input  [3:0]   io_recv_sync,
  input          io_recv_sync_phase2,
  input          io_signal,
  output         io_signal_ack,
  input  [1:0]   io_local_fpga_id,
  output         io_end,
  input  [31:0]  io_packet_size,
  input  [31:0]  io_level,
  input  [31:0]  io_pending_time,
  input  [31:0]  io_pending_parameter,
  input  [1:0]   io_idol_fpga_num
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  collector_clock; // @[bfs_remote.scala 312:25]
  wire  collector_reset; // @[bfs_remote.scala 312:25]
  wire  collector_io_in_ready; // @[bfs_remote.scala 312:25]
  wire  collector_io_in_valid; // @[bfs_remote.scala 312:25]
  wire [511:0] collector_io_in_bits_tdata; // @[bfs_remote.scala 312:25]
  wire [15:0] collector_io_in_bits_tkeep; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_ready; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_valid; // @[bfs_remote.scala 312:25]
  wire [511:0] collector_io_out_bits_tdata; // @[bfs_remote.scala 312:25]
  wire [15:0] collector_io_out_bits_tkeep; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_bits_tlast; // @[bfs_remote.scala 312:25]
  wire  collector_io_flush; // @[bfs_remote.scala 312:25]
  wire  collector_io_empty; // @[bfs_remote.scala 312:25]
  wire  vertex_in_fifo_s_axis_aclk; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[bfs_remote.scala 319:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[bfs_remote.scala 319:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[bfs_remote.scala 319:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 319:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[bfs_remote.scala 319:30]
  wire [31:0] vertex_in_fifo_axis_rd_data_count; // @[bfs_remote.scala 319:30]
  wire  flow_control_unit_clock; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_reset; // @[bfs_remote.scala 385:33]
  wire [511:0] flow_control_unit_io_data; // @[bfs_remote.scala 385:33]
  wire [15:0] flow_control_unit_io_keep; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_handshake; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_handshake_last; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_period; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_pending_valid; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_pending_bits; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_parameter; // @[bfs_remote.scala 385:33]
  wire [1:0] flow_control_unit_io_idol_fpga_num; // @[bfs_remote.scala 385:33]
  reg [31:0] level; // @[bfs_remote.scala 288:22]
  reg [1:0] local_fpga_id; // @[bfs_remote.scala 290:30]
  reg [31:0] packet_size; // @[bfs_remote.scala 292:28]
  reg [31:0] pending_period; // @[bfs_remote.scala 294:31]
  reg [31:0] pending_parameter; // @[bfs_remote.scala 296:34]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[1:0] == 2'h0 & io_xbar_in_bits_tdata[1:0] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] ? 1'h0 : _filtered_keep_0_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[33:32] == 2'h0 & io_xbar_in_bits_tdata[33:32] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] ? 1'h0 : _filtered_keep_1_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[65:64] == 2'h0 & io_xbar_in_bits_tdata[65:64] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] ? 1'h0 : _filtered_keep_2_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[97:96] == 2'h0 & io_xbar_in_bits_tdata[97:96] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] ? 1'h0 : _filtered_keep_3_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[129:128] == 2'h0 & io_xbar_in_bits_tdata[129:128] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] ? 1'h0 : _filtered_keep_4_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[161:160] == 2'h0 & io_xbar_in_bits_tdata[161:160] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] ? 1'h0 : _filtered_keep_5_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[193:192] == 2'h0 & io_xbar_in_bits_tdata[193:192] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] ? 1'h0 : _filtered_keep_6_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[225:224] == 2'h0 & io_xbar_in_bits_tdata[225:224] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] ? 1'h0 : _filtered_keep_7_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[257:256] == 2'h0 & io_xbar_in_bits_tdata[257:256] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] ? 1'h0 : _filtered_keep_8_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[289:288] == 2'h0 & io_xbar_in_bits_tdata[289:288] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] ? 1'h0 : _filtered_keep_9_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[321:320] == 2'h0 & io_xbar_in_bits_tdata[321:320] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] ? 1'h0 : _filtered_keep_10_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[353:352] == 2'h0 & io_xbar_in_bits_tdata[353:352] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] ? 1'h0 : _filtered_keep_11_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[385:384] == 2'h0 & io_xbar_in_bits_tdata[385:384] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] ? 1'h0 : _filtered_keep_12_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[417:416] == 2'h0 & io_xbar_in_bits_tdata[417:416] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] ? 1'h0 : _filtered_keep_13_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[449:448] == 2'h0 & io_xbar_in_bits_tdata[449:448] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] ? 1'h0 : _filtered_keep_14_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[481:480] == 2'h0 & io_xbar_in_bits_tdata[481:480] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] ? 1'h0 : _filtered_keep_15_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[bfs_remote.scala 306:15]
  wire [7:0] collector_io_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[bfs_remote.scala 314:53]
  wire [7:0] collector_io_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[bfs_remote.scala 314:53]
  reg [31:0] vertex_in_fifo_data_count; // @[bfs_remote.scala 320:42]
  wire  _T_1 = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 321:90]
  wire  _T_2 = vertex_in_fifo_s_axis_tvalid & vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 321:49]
  wire  _T_3 = vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 322:44]
  wire  _T_5 = vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 322:88]
  wire [31:0] _vertex_in_fifo_data_count_T_1 = vertex_in_fifo_data_count + 32'h1; // @[bfs_remote.scala 325:60]
  wire [31:0] _vertex_in_fifo_data_count_T_3 = vertex_in_fifo_data_count - 32'h1; // @[bfs_remote.scala 327:60]
  reg [2:0] sync_status; // @[bfs_remote.scala 345:28]
  reg [31:0] stall_time; // @[bfs_remote.scala 346:27]
  wire  _T_13 = sync_status == 3'h6; // @[bfs_remote.scala 348:20]
  wire [31:0] _stall_time_T_1 = stall_time + 32'h1; // @[bfs_remote.scala 349:30]
  wire  _T_21 = sync_status == 3'h1; // @[bfs_remote.scala 357:26]
  wire  _T_29 = sync_status == 3'h3; // @[bfs_remote.scala 363:26]
  wire [2:0] _GEN_4 = sync_status == 3'h4 & io_signal ? 3'h0 : sync_status; // @[bfs_remote.scala 365:58 bfs_remote.scala 366:17 bfs_remote.scala 345:28]
  wire [2:0] _GEN_5 = sync_status == 3'h3 & _T_1 ? 3'h4 : _GEN_4; // @[bfs_remote.scala 363:95 bfs_remote.scala 364:17]
  wire [2:0] _GEN_6 = _T_13 & stall_time == 32'h1e ? 3'h3 : _GEN_5; // @[bfs_remote.scala 361:71 bfs_remote.scala 362:17]
  wire [2:0] _GEN_7 = sync_status == 3'h2 & io_recv_sync_phase2 ? 3'h6 : _GEN_6; // @[bfs_remote.scala 359:73 bfs_remote.scala 360:17]
  wire  need_to_send_sync = _T_21 | _T_29; // @[bfs_remote.scala 372:66]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = need_to_send_sync ? 16'h1 : collector_io_out_bits_tkeep; // @[bfs_remote.scala 376:40]
  wire [3:0] sync_data_level = level[3:0]; // @[bfs_remote.scala 339:23 bfs_remote.scala 342:19]
  wire [31:0] _vertex_in_fifo_io_s_axis_tdata_T = {1'h1,local_fpga_id,sync_data_level,25'h0}; // @[bfs_remote.scala 378:76]
  reg [31:0] send_count; // @[bfs_remote.scala 382:27]
  reg [31:0] pending_time; // @[bfs_remote.scala 383:29]
  reg [31:0] extra_time; // @[bfs_remote.scala 384:27]
  wire [31:0] _io_remote_out_bits_tlast_T_1 = packet_size - 32'h1; // @[bfs_remote.scala 389:59]
  wire  _io_remote_out_bits_tlast_T_2 = send_count == _io_remote_out_bits_tlast_T_1; // @[bfs_remote.scala 389:42]
  wire  _flow_control_unit_io_handshake_T = io_remote_out_valid & io_remote_out_ready; // @[bfs_remote.scala 392:57]
  wire  _T_34 = pending_time == 32'h0; // @[bfs_remote.scala 399:27]
  wire [31:0] _extra_time_T_1 = extra_time + 32'h1; // @[bfs_remote.scala 400:30]
  wire [31:0] _pending_time_T_2 = flow_control_unit_io_pending_bits - extra_time; // @[bfs_remote.scala 406:46]
  wire [31:0] _pending_time_T_5 = pending_time - 32'h1; // @[bfs_remote.scala 408:34]
  wire [31:0] _send_count_T_1 = send_count + 32'h1; // @[bfs_remote.scala 414:32]
  wire  _T_42 = vertex_in_fifo_data_count >= packet_size & send_count == 32'h0; // @[bfs_remote.scala 417:49]
  wire  _T_44 = _T_42 | send_count != 32'h0; // @[bfs_remote.scala 418:3]
  wire  _GEN_17 = _T_34 & vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 420:31 bfs_remote.scala 421:27 bfs_remote.scala 402:23]
  wire  _GEN_18 = _T_34 & io_remote_out_ready; // @[bfs_remote.scala 420:31 bfs_remote.scala 422:39 bfs_remote.scala 403:35]
  axis_data_collector collector ( // @[bfs_remote.scala 312:25]
    .clock(collector_clock),
    .reset(collector_reset),
    .io_in_ready(collector_io_in_ready),
    .io_in_valid(collector_io_in_valid),
    .io_in_bits_tdata(collector_io_in_bits_tdata),
    .io_in_bits_tkeep(collector_io_in_bits_tkeep),
    .io_out_ready(collector_io_out_ready),
    .io_out_valid(collector_io_out_valid),
    .io_out_bits_tdata(collector_io_out_bits_tdata),
    .io_out_bits_tkeep(collector_io_out_bits_tkeep),
    .io_out_bits_tlast(collector_io_out_bits_tlast),
    .io_flush(collector_io_flush),
    .io_empty(collector_io_empty)
  );
  remote_apply_vid_fifo vertex_in_fifo ( // @[bfs_remote.scala 319:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_in_fifo_axis_rd_data_count)
  );
  flow_control flow_control_unit ( // @[bfs_remote.scala 385:33]
    .clock(flow_control_unit_clock),
    .reset(flow_control_unit_reset),
    .io_data(flow_control_unit_io_data),
    .io_keep(flow_control_unit_io_keep),
    .io_handshake(flow_control_unit_io_handshake),
    .io_handshake_last(flow_control_unit_io_handshake_last),
    .io_period(flow_control_unit_io_period),
    .io_pending_valid(flow_control_unit_io_pending_valid),
    .io_pending_bits(flow_control_unit_io_pending_bits),
    .io_parameter(flow_control_unit_io_parameter),
    .io_idol_fpga_num(flow_control_unit_io_idol_fpga_num)
  );
  assign io_xbar_in_ready = collector_io_in_ready; // @[bfs_remote.scala 317:20]
  assign io_remote_out_valid = (_T_44 | sync_status != 3'h0) & _GEN_17; // @[bfs_remote.scala 419:33 bfs_remote.scala 402:23]
  assign io_remote_out_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 387:28]
  assign io_remote_out_bits_tkeep = vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 386:28]
  assign io_remote_out_bits_tlast = send_count == _io_remote_out_bits_tlast_T_1 | vertex_in_fifo_data_count == 32'h1; // @[bfs_remote.scala 389:66]
  assign io_signal_ack = sync_status == 3'h4; // @[bfs_remote.scala 368:32]
  assign io_end = _T_29 & _T_1; // @[bfs_remote.scala 369:50]
  assign collector_clock = clock;
  assign collector_reset = reset;
  assign collector_io_in_valid = io_xbar_in_valid; // @[bfs_remote.scala 313:25]
  assign collector_io_in_bits_tdata = io_xbar_in_bits_tdata; // @[bfs_remote.scala 315:30]
  assign collector_io_in_bits_tkeep = {collector_io_in_bits_tkeep_hi,collector_io_in_bits_tkeep_lo}; // @[bfs_remote.scala 314:53]
  assign collector_io_out_ready = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 379:26]
  assign collector_io_flush = sync_status == 3'h5; // @[bfs_remote.scala 370:37]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[bfs_remote.scala 373:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[bfs_remote.scala 374:39]
  assign vertex_in_fifo_s_axis_tdata = need_to_send_sync ? {{480'd0}, _vertex_in_fifo_io_s_axis_tdata_T} :
    collector_io_out_bits_tdata; // @[bfs_remote.scala 378:40]
  assign vertex_in_fifo_s_axis_tvalid = collector_io_out_valid | need_to_send_sync; // @[bfs_remote.scala 375:63]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[bfs_remote.scala 376:40]
  assign vertex_in_fifo_s_axis_tlast = 1'h1; // @[bfs_remote.scala 377:34]
  assign vertex_in_fifo_m_axis_tready = (_T_44 | sync_status != 3'h0) & _GEN_18; // @[bfs_remote.scala 419:33 bfs_remote.scala 403:35]
  assign flow_control_unit_clock = clock;
  assign flow_control_unit_reset = reset;
  assign flow_control_unit_io_data = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 390:29]
  assign flow_control_unit_io_keep = vertex_in_fifo_m_axis_tkeep[15:0]; // @[bfs_remote.scala 391:29]
  assign flow_control_unit_io_handshake = io_remote_out_valid & io_remote_out_ready; // @[bfs_remote.scala 392:57]
  assign flow_control_unit_io_handshake_last = io_remote_out_bits_tlast; // @[bfs_remote.scala 393:39]
  assign flow_control_unit_io_period = pending_period; // @[bfs_remote.scala 394:31]
  assign flow_control_unit_io_parameter = pending_parameter; // @[bfs_remote.scala 395:34]
  assign flow_control_unit_io_idol_fpga_num = io_idol_fpga_num; // @[bfs_remote.scala 396:38]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 288:22]
      level <= 32'h0; // @[bfs_remote.scala 288:22]
    end else begin
      level <= io_level; // @[bfs_remote.scala 289:9]
    end
    if (reset) begin // @[bfs_remote.scala 290:30]
      local_fpga_id <= 2'h0; // @[bfs_remote.scala 290:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[bfs_remote.scala 291:17]
    end
    if (reset) begin // @[bfs_remote.scala 292:28]
      packet_size <= 32'h0; // @[bfs_remote.scala 292:28]
    end else begin
      packet_size <= io_packet_size; // @[bfs_remote.scala 293:15]
    end
    if (reset) begin // @[bfs_remote.scala 294:31]
      pending_period <= 32'h0; // @[bfs_remote.scala 294:31]
    end else begin
      pending_period <= io_pending_time; // @[bfs_remote.scala 295:18]
    end
    if (reset) begin // @[bfs_remote.scala 296:34]
      pending_parameter <= 32'h0; // @[bfs_remote.scala 296:34]
    end else begin
      pending_parameter <= io_pending_parameter; // @[bfs_remote.scala 297:21]
    end
    if (reset) begin // @[bfs_remote.scala 320:42]
      vertex_in_fifo_data_count <= 32'h0; // @[bfs_remote.scala 320:42]
    end else if (!(_T_2 & vertex_in_fifo_m_axis_tvalid & vertex_in_fifo_m_axis_tready)) begin // @[bfs_remote.scala 322:92]
      if (_T_2) begin // @[bfs_remote.scala 324:99]
        vertex_in_fifo_data_count <= _vertex_in_fifo_data_count_T_1; // @[bfs_remote.scala 325:31]
      end else if (_T_3 & _T_5) begin // @[bfs_remote.scala 326:99]
        vertex_in_fifo_data_count <= _vertex_in_fifo_data_count_T_3; // @[bfs_remote.scala 327:31]
      end
    end
    if (reset) begin // @[bfs_remote.scala 345:28]
      sync_status <= 3'h0; // @[bfs_remote.scala 345:28]
    end else if (sync_status == 3'h0 & &io_recv_sync & local_fpga_id != 2'h0) begin // @[bfs_remote.scala 353:90]
      sync_status <= 3'h5; // @[bfs_remote.scala 354:17]
    end else if (sync_status == 3'h5 & collector_io_empty) begin // @[bfs_remote.scala 355:61]
      sync_status <= 3'h1; // @[bfs_remote.scala 356:17]
    end else if (sync_status == 3'h1 & _T_1) begin // @[bfs_remote.scala 357:95]
      sync_status <= 3'h2; // @[bfs_remote.scala 358:17]
    end else begin
      sync_status <= _GEN_7;
    end
    if (reset) begin // @[bfs_remote.scala 346:27]
      stall_time <= 32'h0; // @[bfs_remote.scala 346:27]
    end else if (sync_status == 3'h6) begin // @[bfs_remote.scala 348:42]
      stall_time <= _stall_time_T_1; // @[bfs_remote.scala 349:16]
    end else begin
      stall_time <= 32'h0; // @[bfs_remote.scala 351:16]
    end
    if (reset) begin // @[bfs_remote.scala 382:27]
      send_count <= 32'h0; // @[bfs_remote.scala 382:27]
    end else if (_flow_control_unit_io_handshake_T) begin // @[bfs_remote.scala 410:51]
      if (_io_remote_out_bits_tlast_T_2) begin // @[bfs_remote.scala 411:45]
        send_count <= 32'h0; // @[bfs_remote.scala 412:18]
      end else begin
        send_count <= _send_count_T_1; // @[bfs_remote.scala 414:18]
      end
    end
    if (reset) begin // @[bfs_remote.scala 383:29]
      pending_time <= 32'h0; // @[bfs_remote.scala 383:29]
    end else if (flow_control_unit_io_pending_valid) begin // @[bfs_remote.scala 404:43]
      if (extra_time > flow_control_unit_io_pending_bits) begin // @[bfs_remote.scala 405:24]
        pending_time <= 32'h0;
      end else begin
        pending_time <= _pending_time_T_2;
      end
    end else if (pending_time != 32'h0) begin // @[bfs_remote.scala 407:35]
      pending_time <= _pending_time_T_5; // @[bfs_remote.scala 408:18]
    end
    if (reset) begin // @[bfs_remote.scala 384:27]
      extra_time <= 32'h0; // @[bfs_remote.scala 384:27]
    end else if (flow_control_unit_io_pending_valid) begin // @[bfs_remote.scala 397:43]
      extra_time <= 32'h0; // @[bfs_remote.scala 398:16]
    end else if (pending_time == 32'h0) begin // @[bfs_remote.scala 399:35]
      extra_time <= _extra_time_T_1; // @[bfs_remote.scala 400:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  level = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  local_fpga_id = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  packet_size = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  pending_period = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pending_parameter = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  vertex_in_fifo_data_count = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  sync_status = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  stall_time = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  send_count = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  pending_time = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  extra_time = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Remote_Apply_1(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_remote_out_ready,
  output         io_remote_out_valid,
  output [511:0] io_remote_out_bits_tdata,
  output [63:0]  io_remote_out_bits_tkeep,
  output         io_remote_out_bits_tlast,
  input  [3:0]   io_recv_sync,
  input          io_recv_sync_phase2,
  input          io_signal,
  output         io_signal_ack,
  input  [1:0]   io_local_fpga_id,
  output         io_end,
  input  [31:0]  io_packet_size,
  input  [31:0]  io_level,
  input  [31:0]  io_pending_time,
  input  [31:0]  io_pending_parameter,
  input  [1:0]   io_idol_fpga_num
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  collector_clock; // @[bfs_remote.scala 312:25]
  wire  collector_reset; // @[bfs_remote.scala 312:25]
  wire  collector_io_in_ready; // @[bfs_remote.scala 312:25]
  wire  collector_io_in_valid; // @[bfs_remote.scala 312:25]
  wire [511:0] collector_io_in_bits_tdata; // @[bfs_remote.scala 312:25]
  wire [15:0] collector_io_in_bits_tkeep; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_ready; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_valid; // @[bfs_remote.scala 312:25]
  wire [511:0] collector_io_out_bits_tdata; // @[bfs_remote.scala 312:25]
  wire [15:0] collector_io_out_bits_tkeep; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_bits_tlast; // @[bfs_remote.scala 312:25]
  wire  collector_io_flush; // @[bfs_remote.scala 312:25]
  wire  collector_io_empty; // @[bfs_remote.scala 312:25]
  wire  vertex_in_fifo_s_axis_aclk; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[bfs_remote.scala 319:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[bfs_remote.scala 319:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[bfs_remote.scala 319:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 319:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[bfs_remote.scala 319:30]
  wire [31:0] vertex_in_fifo_axis_rd_data_count; // @[bfs_remote.scala 319:30]
  wire  flow_control_unit_clock; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_reset; // @[bfs_remote.scala 385:33]
  wire [511:0] flow_control_unit_io_data; // @[bfs_remote.scala 385:33]
  wire [15:0] flow_control_unit_io_keep; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_handshake; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_handshake_last; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_period; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_pending_valid; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_pending_bits; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_parameter; // @[bfs_remote.scala 385:33]
  wire [1:0] flow_control_unit_io_idol_fpga_num; // @[bfs_remote.scala 385:33]
  reg [31:0] level; // @[bfs_remote.scala 288:22]
  reg [1:0] local_fpga_id; // @[bfs_remote.scala 290:30]
  reg [31:0] packet_size; // @[bfs_remote.scala 292:28]
  reg [31:0] pending_period; // @[bfs_remote.scala 294:31]
  reg [31:0] pending_parameter; // @[bfs_remote.scala 296:34]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[1:0] == 2'h1 & io_xbar_in_bits_tdata[1:0] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] ? 1'h0 : _filtered_keep_0_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[33:32] == 2'h1 & io_xbar_in_bits_tdata[33:32] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] ? 1'h0 : _filtered_keep_1_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[65:64] == 2'h1 & io_xbar_in_bits_tdata[65:64] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] ? 1'h0 : _filtered_keep_2_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[97:96] == 2'h1 & io_xbar_in_bits_tdata[97:96] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] ? 1'h0 : _filtered_keep_3_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[129:128] == 2'h1 & io_xbar_in_bits_tdata[129:128] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] ? 1'h0 : _filtered_keep_4_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[161:160] == 2'h1 & io_xbar_in_bits_tdata[161:160] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] ? 1'h0 : _filtered_keep_5_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[193:192] == 2'h1 & io_xbar_in_bits_tdata[193:192] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] ? 1'h0 : _filtered_keep_6_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[225:224] == 2'h1 & io_xbar_in_bits_tdata[225:224] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] ? 1'h0 : _filtered_keep_7_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[257:256] == 2'h1 & io_xbar_in_bits_tdata[257:256] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] ? 1'h0 : _filtered_keep_8_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[289:288] == 2'h1 & io_xbar_in_bits_tdata[289:288] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] ? 1'h0 : _filtered_keep_9_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[321:320] == 2'h1 & io_xbar_in_bits_tdata[321:320] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] ? 1'h0 : _filtered_keep_10_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[353:352] == 2'h1 & io_xbar_in_bits_tdata[353:352] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] ? 1'h0 : _filtered_keep_11_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[385:384] == 2'h1 & io_xbar_in_bits_tdata[385:384] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] ? 1'h0 : _filtered_keep_12_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[417:416] == 2'h1 & io_xbar_in_bits_tdata[417:416] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] ? 1'h0 : _filtered_keep_13_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[449:448] == 2'h1 & io_xbar_in_bits_tdata[449:448] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] ? 1'h0 : _filtered_keep_14_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[481:480] == 2'h1 & io_xbar_in_bits_tdata[481:480] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] ? 1'h0 : _filtered_keep_15_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[bfs_remote.scala 306:15]
  wire [7:0] collector_io_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[bfs_remote.scala 314:53]
  wire [7:0] collector_io_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[bfs_remote.scala 314:53]
  reg [31:0] vertex_in_fifo_data_count; // @[bfs_remote.scala 320:42]
  wire  _T_1 = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 321:90]
  wire  _T_2 = vertex_in_fifo_s_axis_tvalid & vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 321:49]
  wire  _T_3 = vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 322:44]
  wire  _T_5 = vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 322:88]
  wire [31:0] _vertex_in_fifo_data_count_T_1 = vertex_in_fifo_data_count + 32'h1; // @[bfs_remote.scala 325:60]
  wire [31:0] _vertex_in_fifo_data_count_T_3 = vertex_in_fifo_data_count - 32'h1; // @[bfs_remote.scala 327:60]
  reg [2:0] sync_status; // @[bfs_remote.scala 345:28]
  reg [31:0] stall_time; // @[bfs_remote.scala 346:27]
  wire  _T_13 = sync_status == 3'h6; // @[bfs_remote.scala 348:20]
  wire [31:0] _stall_time_T_1 = stall_time + 32'h1; // @[bfs_remote.scala 349:30]
  wire  _T_21 = sync_status == 3'h1; // @[bfs_remote.scala 357:26]
  wire  _T_29 = sync_status == 3'h3; // @[bfs_remote.scala 363:26]
  wire [2:0] _GEN_4 = sync_status == 3'h4 & io_signal ? 3'h0 : sync_status; // @[bfs_remote.scala 365:58 bfs_remote.scala 366:17 bfs_remote.scala 345:28]
  wire [2:0] _GEN_5 = sync_status == 3'h3 & _T_1 ? 3'h4 : _GEN_4; // @[bfs_remote.scala 363:95 bfs_remote.scala 364:17]
  wire [2:0] _GEN_6 = _T_13 & stall_time == 32'h1e ? 3'h3 : _GEN_5; // @[bfs_remote.scala 361:71 bfs_remote.scala 362:17]
  wire [2:0] _GEN_7 = sync_status == 3'h2 & io_recv_sync_phase2 ? 3'h6 : _GEN_6; // @[bfs_remote.scala 359:73 bfs_remote.scala 360:17]
  wire  need_to_send_sync = _T_21 | _T_29; // @[bfs_remote.scala 372:66]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = need_to_send_sync ? 16'h1 : collector_io_out_bits_tkeep; // @[bfs_remote.scala 376:40]
  wire [3:0] sync_data_level = level[3:0]; // @[bfs_remote.scala 339:23 bfs_remote.scala 342:19]
  wire [31:0] _vertex_in_fifo_io_s_axis_tdata_T = {1'h1,local_fpga_id,sync_data_level,25'h0}; // @[bfs_remote.scala 378:76]
  reg [31:0] send_count; // @[bfs_remote.scala 382:27]
  reg [31:0] pending_time; // @[bfs_remote.scala 383:29]
  reg [31:0] extra_time; // @[bfs_remote.scala 384:27]
  wire [31:0] _io_remote_out_bits_tlast_T_1 = packet_size - 32'h1; // @[bfs_remote.scala 389:59]
  wire  _io_remote_out_bits_tlast_T_2 = send_count == _io_remote_out_bits_tlast_T_1; // @[bfs_remote.scala 389:42]
  wire  _flow_control_unit_io_handshake_T = io_remote_out_valid & io_remote_out_ready; // @[bfs_remote.scala 392:57]
  wire  _T_34 = pending_time == 32'h0; // @[bfs_remote.scala 399:27]
  wire [31:0] _extra_time_T_1 = extra_time + 32'h1; // @[bfs_remote.scala 400:30]
  wire [31:0] _pending_time_T_2 = flow_control_unit_io_pending_bits - extra_time; // @[bfs_remote.scala 406:46]
  wire [31:0] _pending_time_T_5 = pending_time - 32'h1; // @[bfs_remote.scala 408:34]
  wire [31:0] _send_count_T_1 = send_count + 32'h1; // @[bfs_remote.scala 414:32]
  wire  _T_42 = vertex_in_fifo_data_count >= packet_size & send_count == 32'h0; // @[bfs_remote.scala 417:49]
  wire  _T_44 = _T_42 | send_count != 32'h0; // @[bfs_remote.scala 418:3]
  wire  _GEN_17 = _T_34 & vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 420:31 bfs_remote.scala 421:27 bfs_remote.scala 402:23]
  wire  _GEN_18 = _T_34 & io_remote_out_ready; // @[bfs_remote.scala 420:31 bfs_remote.scala 422:39 bfs_remote.scala 403:35]
  axis_data_collector collector ( // @[bfs_remote.scala 312:25]
    .clock(collector_clock),
    .reset(collector_reset),
    .io_in_ready(collector_io_in_ready),
    .io_in_valid(collector_io_in_valid),
    .io_in_bits_tdata(collector_io_in_bits_tdata),
    .io_in_bits_tkeep(collector_io_in_bits_tkeep),
    .io_out_ready(collector_io_out_ready),
    .io_out_valid(collector_io_out_valid),
    .io_out_bits_tdata(collector_io_out_bits_tdata),
    .io_out_bits_tkeep(collector_io_out_bits_tkeep),
    .io_out_bits_tlast(collector_io_out_bits_tlast),
    .io_flush(collector_io_flush),
    .io_empty(collector_io_empty)
  );
  remote_apply_vid_fifo vertex_in_fifo ( // @[bfs_remote.scala 319:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_in_fifo_axis_rd_data_count)
  );
  flow_control flow_control_unit ( // @[bfs_remote.scala 385:33]
    .clock(flow_control_unit_clock),
    .reset(flow_control_unit_reset),
    .io_data(flow_control_unit_io_data),
    .io_keep(flow_control_unit_io_keep),
    .io_handshake(flow_control_unit_io_handshake),
    .io_handshake_last(flow_control_unit_io_handshake_last),
    .io_period(flow_control_unit_io_period),
    .io_pending_valid(flow_control_unit_io_pending_valid),
    .io_pending_bits(flow_control_unit_io_pending_bits),
    .io_parameter(flow_control_unit_io_parameter),
    .io_idol_fpga_num(flow_control_unit_io_idol_fpga_num)
  );
  assign io_xbar_in_ready = collector_io_in_ready; // @[bfs_remote.scala 317:20]
  assign io_remote_out_valid = (_T_44 | sync_status != 3'h0) & _GEN_17; // @[bfs_remote.scala 419:33 bfs_remote.scala 402:23]
  assign io_remote_out_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 387:28]
  assign io_remote_out_bits_tkeep = vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 386:28]
  assign io_remote_out_bits_tlast = send_count == _io_remote_out_bits_tlast_T_1 | vertex_in_fifo_data_count == 32'h1; // @[bfs_remote.scala 389:66]
  assign io_signal_ack = sync_status == 3'h4; // @[bfs_remote.scala 368:32]
  assign io_end = _T_29 & _T_1; // @[bfs_remote.scala 369:50]
  assign collector_clock = clock;
  assign collector_reset = reset;
  assign collector_io_in_valid = io_xbar_in_valid; // @[bfs_remote.scala 313:25]
  assign collector_io_in_bits_tdata = io_xbar_in_bits_tdata; // @[bfs_remote.scala 315:30]
  assign collector_io_in_bits_tkeep = {collector_io_in_bits_tkeep_hi,collector_io_in_bits_tkeep_lo}; // @[bfs_remote.scala 314:53]
  assign collector_io_out_ready = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 379:26]
  assign collector_io_flush = sync_status == 3'h5; // @[bfs_remote.scala 370:37]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[bfs_remote.scala 373:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[bfs_remote.scala 374:39]
  assign vertex_in_fifo_s_axis_tdata = need_to_send_sync ? {{480'd0}, _vertex_in_fifo_io_s_axis_tdata_T} :
    collector_io_out_bits_tdata; // @[bfs_remote.scala 378:40]
  assign vertex_in_fifo_s_axis_tvalid = collector_io_out_valid | need_to_send_sync; // @[bfs_remote.scala 375:63]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[bfs_remote.scala 376:40]
  assign vertex_in_fifo_s_axis_tlast = 1'h1; // @[bfs_remote.scala 377:34]
  assign vertex_in_fifo_m_axis_tready = (_T_44 | sync_status != 3'h0) & _GEN_18; // @[bfs_remote.scala 419:33 bfs_remote.scala 403:35]
  assign flow_control_unit_clock = clock;
  assign flow_control_unit_reset = reset;
  assign flow_control_unit_io_data = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 390:29]
  assign flow_control_unit_io_keep = vertex_in_fifo_m_axis_tkeep[15:0]; // @[bfs_remote.scala 391:29]
  assign flow_control_unit_io_handshake = io_remote_out_valid & io_remote_out_ready; // @[bfs_remote.scala 392:57]
  assign flow_control_unit_io_handshake_last = io_remote_out_bits_tlast; // @[bfs_remote.scala 393:39]
  assign flow_control_unit_io_period = pending_period; // @[bfs_remote.scala 394:31]
  assign flow_control_unit_io_parameter = pending_parameter; // @[bfs_remote.scala 395:34]
  assign flow_control_unit_io_idol_fpga_num = io_idol_fpga_num; // @[bfs_remote.scala 396:38]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 288:22]
      level <= 32'h0; // @[bfs_remote.scala 288:22]
    end else begin
      level <= io_level; // @[bfs_remote.scala 289:9]
    end
    if (reset) begin // @[bfs_remote.scala 290:30]
      local_fpga_id <= 2'h0; // @[bfs_remote.scala 290:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[bfs_remote.scala 291:17]
    end
    if (reset) begin // @[bfs_remote.scala 292:28]
      packet_size <= 32'h0; // @[bfs_remote.scala 292:28]
    end else begin
      packet_size <= io_packet_size; // @[bfs_remote.scala 293:15]
    end
    if (reset) begin // @[bfs_remote.scala 294:31]
      pending_period <= 32'h0; // @[bfs_remote.scala 294:31]
    end else begin
      pending_period <= io_pending_time; // @[bfs_remote.scala 295:18]
    end
    if (reset) begin // @[bfs_remote.scala 296:34]
      pending_parameter <= 32'h0; // @[bfs_remote.scala 296:34]
    end else begin
      pending_parameter <= io_pending_parameter; // @[bfs_remote.scala 297:21]
    end
    if (reset) begin // @[bfs_remote.scala 320:42]
      vertex_in_fifo_data_count <= 32'h0; // @[bfs_remote.scala 320:42]
    end else if (!(_T_2 & vertex_in_fifo_m_axis_tvalid & vertex_in_fifo_m_axis_tready)) begin // @[bfs_remote.scala 322:92]
      if (_T_2) begin // @[bfs_remote.scala 324:99]
        vertex_in_fifo_data_count <= _vertex_in_fifo_data_count_T_1; // @[bfs_remote.scala 325:31]
      end else if (_T_3 & _T_5) begin // @[bfs_remote.scala 326:99]
        vertex_in_fifo_data_count <= _vertex_in_fifo_data_count_T_3; // @[bfs_remote.scala 327:31]
      end
    end
    if (reset) begin // @[bfs_remote.scala 345:28]
      sync_status <= 3'h0; // @[bfs_remote.scala 345:28]
    end else if (sync_status == 3'h0 & &io_recv_sync & local_fpga_id != 2'h1) begin // @[bfs_remote.scala 353:90]
      sync_status <= 3'h5; // @[bfs_remote.scala 354:17]
    end else if (sync_status == 3'h5 & collector_io_empty) begin // @[bfs_remote.scala 355:61]
      sync_status <= 3'h1; // @[bfs_remote.scala 356:17]
    end else if (sync_status == 3'h1 & _T_1) begin // @[bfs_remote.scala 357:95]
      sync_status <= 3'h2; // @[bfs_remote.scala 358:17]
    end else begin
      sync_status <= _GEN_7;
    end
    if (reset) begin // @[bfs_remote.scala 346:27]
      stall_time <= 32'h0; // @[bfs_remote.scala 346:27]
    end else if (sync_status == 3'h6) begin // @[bfs_remote.scala 348:42]
      stall_time <= _stall_time_T_1; // @[bfs_remote.scala 349:16]
    end else begin
      stall_time <= 32'h0; // @[bfs_remote.scala 351:16]
    end
    if (reset) begin // @[bfs_remote.scala 382:27]
      send_count <= 32'h0; // @[bfs_remote.scala 382:27]
    end else if (_flow_control_unit_io_handshake_T) begin // @[bfs_remote.scala 410:51]
      if (_io_remote_out_bits_tlast_T_2) begin // @[bfs_remote.scala 411:45]
        send_count <= 32'h0; // @[bfs_remote.scala 412:18]
      end else begin
        send_count <= _send_count_T_1; // @[bfs_remote.scala 414:18]
      end
    end
    if (reset) begin // @[bfs_remote.scala 383:29]
      pending_time <= 32'h0; // @[bfs_remote.scala 383:29]
    end else if (flow_control_unit_io_pending_valid) begin // @[bfs_remote.scala 404:43]
      if (extra_time > flow_control_unit_io_pending_bits) begin // @[bfs_remote.scala 405:24]
        pending_time <= 32'h0;
      end else begin
        pending_time <= _pending_time_T_2;
      end
    end else if (pending_time != 32'h0) begin // @[bfs_remote.scala 407:35]
      pending_time <= _pending_time_T_5; // @[bfs_remote.scala 408:18]
    end
    if (reset) begin // @[bfs_remote.scala 384:27]
      extra_time <= 32'h0; // @[bfs_remote.scala 384:27]
    end else if (flow_control_unit_io_pending_valid) begin // @[bfs_remote.scala 397:43]
      extra_time <= 32'h0; // @[bfs_remote.scala 398:16]
    end else if (pending_time == 32'h0) begin // @[bfs_remote.scala 399:35]
      extra_time <= _extra_time_T_1; // @[bfs_remote.scala 400:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  level = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  local_fpga_id = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  packet_size = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  pending_period = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pending_parameter = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  vertex_in_fifo_data_count = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  sync_status = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  stall_time = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  send_count = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  pending_time = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  extra_time = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Remote_Apply_2(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_remote_out_ready,
  output         io_remote_out_valid,
  output [511:0] io_remote_out_bits_tdata,
  output [63:0]  io_remote_out_bits_tkeep,
  output         io_remote_out_bits_tlast,
  input  [3:0]   io_recv_sync,
  input          io_recv_sync_phase2,
  input          io_signal,
  output         io_signal_ack,
  input  [1:0]   io_local_fpga_id,
  output         io_end,
  input  [31:0]  io_packet_size,
  input  [31:0]  io_level,
  input  [31:0]  io_pending_time,
  input  [31:0]  io_pending_parameter,
  input  [1:0]   io_idol_fpga_num
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  collector_clock; // @[bfs_remote.scala 312:25]
  wire  collector_reset; // @[bfs_remote.scala 312:25]
  wire  collector_io_in_ready; // @[bfs_remote.scala 312:25]
  wire  collector_io_in_valid; // @[bfs_remote.scala 312:25]
  wire [511:0] collector_io_in_bits_tdata; // @[bfs_remote.scala 312:25]
  wire [15:0] collector_io_in_bits_tkeep; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_ready; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_valid; // @[bfs_remote.scala 312:25]
  wire [511:0] collector_io_out_bits_tdata; // @[bfs_remote.scala 312:25]
  wire [15:0] collector_io_out_bits_tkeep; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_bits_tlast; // @[bfs_remote.scala 312:25]
  wire  collector_io_flush; // @[bfs_remote.scala 312:25]
  wire  collector_io_empty; // @[bfs_remote.scala 312:25]
  wire  vertex_in_fifo_s_axis_aclk; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[bfs_remote.scala 319:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[bfs_remote.scala 319:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[bfs_remote.scala 319:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 319:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[bfs_remote.scala 319:30]
  wire [31:0] vertex_in_fifo_axis_rd_data_count; // @[bfs_remote.scala 319:30]
  wire  flow_control_unit_clock; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_reset; // @[bfs_remote.scala 385:33]
  wire [511:0] flow_control_unit_io_data; // @[bfs_remote.scala 385:33]
  wire [15:0] flow_control_unit_io_keep; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_handshake; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_handshake_last; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_period; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_pending_valid; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_pending_bits; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_parameter; // @[bfs_remote.scala 385:33]
  wire [1:0] flow_control_unit_io_idol_fpga_num; // @[bfs_remote.scala 385:33]
  reg [31:0] level; // @[bfs_remote.scala 288:22]
  reg [1:0] local_fpga_id; // @[bfs_remote.scala 290:30]
  reg [31:0] packet_size; // @[bfs_remote.scala 292:28]
  reg [31:0] pending_period; // @[bfs_remote.scala 294:31]
  reg [31:0] pending_parameter; // @[bfs_remote.scala 296:34]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[1:0] == 2'h2 & io_xbar_in_bits_tdata[1:0] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] ? 1'h0 : _filtered_keep_0_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[33:32] == 2'h2 & io_xbar_in_bits_tdata[33:32] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] ? 1'h0 : _filtered_keep_1_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[65:64] == 2'h2 & io_xbar_in_bits_tdata[65:64] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] ? 1'h0 : _filtered_keep_2_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[97:96] == 2'h2 & io_xbar_in_bits_tdata[97:96] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] ? 1'h0 : _filtered_keep_3_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[129:128] == 2'h2 & io_xbar_in_bits_tdata[129:128] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] ? 1'h0 : _filtered_keep_4_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[161:160] == 2'h2 & io_xbar_in_bits_tdata[161:160] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] ? 1'h0 : _filtered_keep_5_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[193:192] == 2'h2 & io_xbar_in_bits_tdata[193:192] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] ? 1'h0 : _filtered_keep_6_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[225:224] == 2'h2 & io_xbar_in_bits_tdata[225:224] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] ? 1'h0 : _filtered_keep_7_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[257:256] == 2'h2 & io_xbar_in_bits_tdata[257:256] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] ? 1'h0 : _filtered_keep_8_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[289:288] == 2'h2 & io_xbar_in_bits_tdata[289:288] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] ? 1'h0 : _filtered_keep_9_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[321:320] == 2'h2 & io_xbar_in_bits_tdata[321:320] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] ? 1'h0 : _filtered_keep_10_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[353:352] == 2'h2 & io_xbar_in_bits_tdata[353:352] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] ? 1'h0 : _filtered_keep_11_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[385:384] == 2'h2 & io_xbar_in_bits_tdata[385:384] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] ? 1'h0 : _filtered_keep_12_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[417:416] == 2'h2 & io_xbar_in_bits_tdata[417:416] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] ? 1'h0 : _filtered_keep_13_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[449:448] == 2'h2 & io_xbar_in_bits_tdata[449:448] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] ? 1'h0 : _filtered_keep_14_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[481:480] == 2'h2 & io_xbar_in_bits_tdata[481:480] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] ? 1'h0 : _filtered_keep_15_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[bfs_remote.scala 306:15]
  wire [7:0] collector_io_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[bfs_remote.scala 314:53]
  wire [7:0] collector_io_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[bfs_remote.scala 314:53]
  reg [31:0] vertex_in_fifo_data_count; // @[bfs_remote.scala 320:42]
  wire  _T_1 = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 321:90]
  wire  _T_2 = vertex_in_fifo_s_axis_tvalid & vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 321:49]
  wire  _T_3 = vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 322:44]
  wire  _T_5 = vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 322:88]
  wire [31:0] _vertex_in_fifo_data_count_T_1 = vertex_in_fifo_data_count + 32'h1; // @[bfs_remote.scala 325:60]
  wire [31:0] _vertex_in_fifo_data_count_T_3 = vertex_in_fifo_data_count - 32'h1; // @[bfs_remote.scala 327:60]
  reg [2:0] sync_status; // @[bfs_remote.scala 345:28]
  reg [31:0] stall_time; // @[bfs_remote.scala 346:27]
  wire  _T_13 = sync_status == 3'h6; // @[bfs_remote.scala 348:20]
  wire [31:0] _stall_time_T_1 = stall_time + 32'h1; // @[bfs_remote.scala 349:30]
  wire  _T_21 = sync_status == 3'h1; // @[bfs_remote.scala 357:26]
  wire  _T_29 = sync_status == 3'h3; // @[bfs_remote.scala 363:26]
  wire [2:0] _GEN_4 = sync_status == 3'h4 & io_signal ? 3'h0 : sync_status; // @[bfs_remote.scala 365:58 bfs_remote.scala 366:17 bfs_remote.scala 345:28]
  wire [2:0] _GEN_5 = sync_status == 3'h3 & _T_1 ? 3'h4 : _GEN_4; // @[bfs_remote.scala 363:95 bfs_remote.scala 364:17]
  wire [2:0] _GEN_6 = _T_13 & stall_time == 32'h1e ? 3'h3 : _GEN_5; // @[bfs_remote.scala 361:71 bfs_remote.scala 362:17]
  wire [2:0] _GEN_7 = sync_status == 3'h2 & io_recv_sync_phase2 ? 3'h6 : _GEN_6; // @[bfs_remote.scala 359:73 bfs_remote.scala 360:17]
  wire  need_to_send_sync = _T_21 | _T_29; // @[bfs_remote.scala 372:66]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = need_to_send_sync ? 16'h1 : collector_io_out_bits_tkeep; // @[bfs_remote.scala 376:40]
  wire [3:0] sync_data_level = level[3:0]; // @[bfs_remote.scala 339:23 bfs_remote.scala 342:19]
  wire [31:0] _vertex_in_fifo_io_s_axis_tdata_T = {1'h1,local_fpga_id,sync_data_level,25'h0}; // @[bfs_remote.scala 378:76]
  reg [31:0] send_count; // @[bfs_remote.scala 382:27]
  reg [31:0] pending_time; // @[bfs_remote.scala 383:29]
  reg [31:0] extra_time; // @[bfs_remote.scala 384:27]
  wire [31:0] _io_remote_out_bits_tlast_T_1 = packet_size - 32'h1; // @[bfs_remote.scala 389:59]
  wire  _io_remote_out_bits_tlast_T_2 = send_count == _io_remote_out_bits_tlast_T_1; // @[bfs_remote.scala 389:42]
  wire  _flow_control_unit_io_handshake_T = io_remote_out_valid & io_remote_out_ready; // @[bfs_remote.scala 392:57]
  wire  _T_34 = pending_time == 32'h0; // @[bfs_remote.scala 399:27]
  wire [31:0] _extra_time_T_1 = extra_time + 32'h1; // @[bfs_remote.scala 400:30]
  wire [31:0] _pending_time_T_2 = flow_control_unit_io_pending_bits - extra_time; // @[bfs_remote.scala 406:46]
  wire [31:0] _pending_time_T_5 = pending_time - 32'h1; // @[bfs_remote.scala 408:34]
  wire [31:0] _send_count_T_1 = send_count + 32'h1; // @[bfs_remote.scala 414:32]
  wire  _T_42 = vertex_in_fifo_data_count >= packet_size & send_count == 32'h0; // @[bfs_remote.scala 417:49]
  wire  _T_44 = _T_42 | send_count != 32'h0; // @[bfs_remote.scala 418:3]
  wire  _GEN_17 = _T_34 & vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 420:31 bfs_remote.scala 421:27 bfs_remote.scala 402:23]
  wire  _GEN_18 = _T_34 & io_remote_out_ready; // @[bfs_remote.scala 420:31 bfs_remote.scala 422:39 bfs_remote.scala 403:35]
  axis_data_collector collector ( // @[bfs_remote.scala 312:25]
    .clock(collector_clock),
    .reset(collector_reset),
    .io_in_ready(collector_io_in_ready),
    .io_in_valid(collector_io_in_valid),
    .io_in_bits_tdata(collector_io_in_bits_tdata),
    .io_in_bits_tkeep(collector_io_in_bits_tkeep),
    .io_out_ready(collector_io_out_ready),
    .io_out_valid(collector_io_out_valid),
    .io_out_bits_tdata(collector_io_out_bits_tdata),
    .io_out_bits_tkeep(collector_io_out_bits_tkeep),
    .io_out_bits_tlast(collector_io_out_bits_tlast),
    .io_flush(collector_io_flush),
    .io_empty(collector_io_empty)
  );
  remote_apply_vid_fifo vertex_in_fifo ( // @[bfs_remote.scala 319:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_in_fifo_axis_rd_data_count)
  );
  flow_control flow_control_unit ( // @[bfs_remote.scala 385:33]
    .clock(flow_control_unit_clock),
    .reset(flow_control_unit_reset),
    .io_data(flow_control_unit_io_data),
    .io_keep(flow_control_unit_io_keep),
    .io_handshake(flow_control_unit_io_handshake),
    .io_handshake_last(flow_control_unit_io_handshake_last),
    .io_period(flow_control_unit_io_period),
    .io_pending_valid(flow_control_unit_io_pending_valid),
    .io_pending_bits(flow_control_unit_io_pending_bits),
    .io_parameter(flow_control_unit_io_parameter),
    .io_idol_fpga_num(flow_control_unit_io_idol_fpga_num)
  );
  assign io_xbar_in_ready = collector_io_in_ready; // @[bfs_remote.scala 317:20]
  assign io_remote_out_valid = (_T_44 | sync_status != 3'h0) & _GEN_17; // @[bfs_remote.scala 419:33 bfs_remote.scala 402:23]
  assign io_remote_out_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 387:28]
  assign io_remote_out_bits_tkeep = vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 386:28]
  assign io_remote_out_bits_tlast = send_count == _io_remote_out_bits_tlast_T_1 | vertex_in_fifo_data_count == 32'h1; // @[bfs_remote.scala 389:66]
  assign io_signal_ack = sync_status == 3'h4; // @[bfs_remote.scala 368:32]
  assign io_end = _T_29 & _T_1; // @[bfs_remote.scala 369:50]
  assign collector_clock = clock;
  assign collector_reset = reset;
  assign collector_io_in_valid = io_xbar_in_valid; // @[bfs_remote.scala 313:25]
  assign collector_io_in_bits_tdata = io_xbar_in_bits_tdata; // @[bfs_remote.scala 315:30]
  assign collector_io_in_bits_tkeep = {collector_io_in_bits_tkeep_hi,collector_io_in_bits_tkeep_lo}; // @[bfs_remote.scala 314:53]
  assign collector_io_out_ready = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 379:26]
  assign collector_io_flush = sync_status == 3'h5; // @[bfs_remote.scala 370:37]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[bfs_remote.scala 373:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[bfs_remote.scala 374:39]
  assign vertex_in_fifo_s_axis_tdata = need_to_send_sync ? {{480'd0}, _vertex_in_fifo_io_s_axis_tdata_T} :
    collector_io_out_bits_tdata; // @[bfs_remote.scala 378:40]
  assign vertex_in_fifo_s_axis_tvalid = collector_io_out_valid | need_to_send_sync; // @[bfs_remote.scala 375:63]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[bfs_remote.scala 376:40]
  assign vertex_in_fifo_s_axis_tlast = 1'h1; // @[bfs_remote.scala 377:34]
  assign vertex_in_fifo_m_axis_tready = (_T_44 | sync_status != 3'h0) & _GEN_18; // @[bfs_remote.scala 419:33 bfs_remote.scala 403:35]
  assign flow_control_unit_clock = clock;
  assign flow_control_unit_reset = reset;
  assign flow_control_unit_io_data = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 390:29]
  assign flow_control_unit_io_keep = vertex_in_fifo_m_axis_tkeep[15:0]; // @[bfs_remote.scala 391:29]
  assign flow_control_unit_io_handshake = io_remote_out_valid & io_remote_out_ready; // @[bfs_remote.scala 392:57]
  assign flow_control_unit_io_handshake_last = io_remote_out_bits_tlast; // @[bfs_remote.scala 393:39]
  assign flow_control_unit_io_period = pending_period; // @[bfs_remote.scala 394:31]
  assign flow_control_unit_io_parameter = pending_parameter; // @[bfs_remote.scala 395:34]
  assign flow_control_unit_io_idol_fpga_num = io_idol_fpga_num; // @[bfs_remote.scala 396:38]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 288:22]
      level <= 32'h0; // @[bfs_remote.scala 288:22]
    end else begin
      level <= io_level; // @[bfs_remote.scala 289:9]
    end
    if (reset) begin // @[bfs_remote.scala 290:30]
      local_fpga_id <= 2'h0; // @[bfs_remote.scala 290:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[bfs_remote.scala 291:17]
    end
    if (reset) begin // @[bfs_remote.scala 292:28]
      packet_size <= 32'h0; // @[bfs_remote.scala 292:28]
    end else begin
      packet_size <= io_packet_size; // @[bfs_remote.scala 293:15]
    end
    if (reset) begin // @[bfs_remote.scala 294:31]
      pending_period <= 32'h0; // @[bfs_remote.scala 294:31]
    end else begin
      pending_period <= io_pending_time; // @[bfs_remote.scala 295:18]
    end
    if (reset) begin // @[bfs_remote.scala 296:34]
      pending_parameter <= 32'h0; // @[bfs_remote.scala 296:34]
    end else begin
      pending_parameter <= io_pending_parameter; // @[bfs_remote.scala 297:21]
    end
    if (reset) begin // @[bfs_remote.scala 320:42]
      vertex_in_fifo_data_count <= 32'h0; // @[bfs_remote.scala 320:42]
    end else if (!(_T_2 & vertex_in_fifo_m_axis_tvalid & vertex_in_fifo_m_axis_tready)) begin // @[bfs_remote.scala 322:92]
      if (_T_2) begin // @[bfs_remote.scala 324:99]
        vertex_in_fifo_data_count <= _vertex_in_fifo_data_count_T_1; // @[bfs_remote.scala 325:31]
      end else if (_T_3 & _T_5) begin // @[bfs_remote.scala 326:99]
        vertex_in_fifo_data_count <= _vertex_in_fifo_data_count_T_3; // @[bfs_remote.scala 327:31]
      end
    end
    if (reset) begin // @[bfs_remote.scala 345:28]
      sync_status <= 3'h0; // @[bfs_remote.scala 345:28]
    end else if (sync_status == 3'h0 & &io_recv_sync & local_fpga_id != 2'h2) begin // @[bfs_remote.scala 353:90]
      sync_status <= 3'h5; // @[bfs_remote.scala 354:17]
    end else if (sync_status == 3'h5 & collector_io_empty) begin // @[bfs_remote.scala 355:61]
      sync_status <= 3'h1; // @[bfs_remote.scala 356:17]
    end else if (sync_status == 3'h1 & _T_1) begin // @[bfs_remote.scala 357:95]
      sync_status <= 3'h2; // @[bfs_remote.scala 358:17]
    end else begin
      sync_status <= _GEN_7;
    end
    if (reset) begin // @[bfs_remote.scala 346:27]
      stall_time <= 32'h0; // @[bfs_remote.scala 346:27]
    end else if (sync_status == 3'h6) begin // @[bfs_remote.scala 348:42]
      stall_time <= _stall_time_T_1; // @[bfs_remote.scala 349:16]
    end else begin
      stall_time <= 32'h0; // @[bfs_remote.scala 351:16]
    end
    if (reset) begin // @[bfs_remote.scala 382:27]
      send_count <= 32'h0; // @[bfs_remote.scala 382:27]
    end else if (_flow_control_unit_io_handshake_T) begin // @[bfs_remote.scala 410:51]
      if (_io_remote_out_bits_tlast_T_2) begin // @[bfs_remote.scala 411:45]
        send_count <= 32'h0; // @[bfs_remote.scala 412:18]
      end else begin
        send_count <= _send_count_T_1; // @[bfs_remote.scala 414:18]
      end
    end
    if (reset) begin // @[bfs_remote.scala 383:29]
      pending_time <= 32'h0; // @[bfs_remote.scala 383:29]
    end else if (flow_control_unit_io_pending_valid) begin // @[bfs_remote.scala 404:43]
      if (extra_time > flow_control_unit_io_pending_bits) begin // @[bfs_remote.scala 405:24]
        pending_time <= 32'h0;
      end else begin
        pending_time <= _pending_time_T_2;
      end
    end else if (pending_time != 32'h0) begin // @[bfs_remote.scala 407:35]
      pending_time <= _pending_time_T_5; // @[bfs_remote.scala 408:18]
    end
    if (reset) begin // @[bfs_remote.scala 384:27]
      extra_time <= 32'h0; // @[bfs_remote.scala 384:27]
    end else if (flow_control_unit_io_pending_valid) begin // @[bfs_remote.scala 397:43]
      extra_time <= 32'h0; // @[bfs_remote.scala 398:16]
    end else if (pending_time == 32'h0) begin // @[bfs_remote.scala 399:35]
      extra_time <= _extra_time_T_1; // @[bfs_remote.scala 400:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  level = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  local_fpga_id = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  packet_size = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  pending_period = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pending_parameter = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  vertex_in_fifo_data_count = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  sync_status = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  stall_time = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  send_count = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  pending_time = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  extra_time = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Remote_Apply_3(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_remote_out_ready,
  output         io_remote_out_valid,
  output [511:0] io_remote_out_bits_tdata,
  output [63:0]  io_remote_out_bits_tkeep,
  output         io_remote_out_bits_tlast,
  input  [3:0]   io_recv_sync,
  input          io_recv_sync_phase2,
  input          io_signal,
  output         io_signal_ack,
  input  [1:0]   io_local_fpga_id,
  output         io_end,
  input  [31:0]  io_packet_size,
  input  [31:0]  io_level,
  input  [31:0]  io_pending_time,
  input  [31:0]  io_pending_parameter,
  input  [1:0]   io_idol_fpga_num
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  collector_clock; // @[bfs_remote.scala 312:25]
  wire  collector_reset; // @[bfs_remote.scala 312:25]
  wire  collector_io_in_ready; // @[bfs_remote.scala 312:25]
  wire  collector_io_in_valid; // @[bfs_remote.scala 312:25]
  wire [511:0] collector_io_in_bits_tdata; // @[bfs_remote.scala 312:25]
  wire [15:0] collector_io_in_bits_tkeep; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_ready; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_valid; // @[bfs_remote.scala 312:25]
  wire [511:0] collector_io_out_bits_tdata; // @[bfs_remote.scala 312:25]
  wire [15:0] collector_io_out_bits_tkeep; // @[bfs_remote.scala 312:25]
  wire  collector_io_out_bits_tlast; // @[bfs_remote.scala 312:25]
  wire  collector_io_flush; // @[bfs_remote.scala 312:25]
  wire  collector_io_empty; // @[bfs_remote.scala 312:25]
  wire  vertex_in_fifo_s_axis_aclk; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[bfs_remote.scala 319:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[bfs_remote.scala 319:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[bfs_remote.scala 319:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 319:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 319:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[bfs_remote.scala 319:30]
  wire [31:0] vertex_in_fifo_axis_rd_data_count; // @[bfs_remote.scala 319:30]
  wire  flow_control_unit_clock; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_reset; // @[bfs_remote.scala 385:33]
  wire [511:0] flow_control_unit_io_data; // @[bfs_remote.scala 385:33]
  wire [15:0] flow_control_unit_io_keep; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_handshake; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_handshake_last; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_period; // @[bfs_remote.scala 385:33]
  wire  flow_control_unit_io_pending_valid; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_pending_bits; // @[bfs_remote.scala 385:33]
  wire [31:0] flow_control_unit_io_parameter; // @[bfs_remote.scala 385:33]
  wire [1:0] flow_control_unit_io_idol_fpga_num; // @[bfs_remote.scala 385:33]
  reg [31:0] level; // @[bfs_remote.scala 288:22]
  reg [1:0] local_fpga_id; // @[bfs_remote.scala 290:30]
  reg [31:0] packet_size; // @[bfs_remote.scala 292:28]
  reg [31:0] pending_period; // @[bfs_remote.scala 294:31]
  reg [31:0] pending_parameter; // @[bfs_remote.scala 296:34]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[1:0] == 2'h3 & io_xbar_in_bits_tdata[1:0] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] ? 1'h0 : _filtered_keep_0_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[33:32] == 2'h3 & io_xbar_in_bits_tdata[33:32] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] ? 1'h0 : _filtered_keep_1_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[65:64] == 2'h3 & io_xbar_in_bits_tdata[65:64] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] ? 1'h0 : _filtered_keep_2_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[97:96] == 2'h3 & io_xbar_in_bits_tdata[97:96] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] ? 1'h0 : _filtered_keep_3_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[129:128] == 2'h3 & io_xbar_in_bits_tdata[129:128] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] ? 1'h0 : _filtered_keep_4_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[161:160] == 2'h3 & io_xbar_in_bits_tdata[161:160] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] ? 1'h0 : _filtered_keep_5_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[193:192] == 2'h3 & io_xbar_in_bits_tdata[193:192] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] ? 1'h0 : _filtered_keep_6_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[225:224] == 2'h3 & io_xbar_in_bits_tdata[225:224] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] ? 1'h0 : _filtered_keep_7_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[257:256] == 2'h3 & io_xbar_in_bits_tdata[257:256] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] ? 1'h0 : _filtered_keep_8_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[289:288] == 2'h3 & io_xbar_in_bits_tdata[289:288] != local_fpga_id; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] ? 1'h0 : _filtered_keep_9_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[321:320] == 2'h3 & io_xbar_in_bits_tdata[321:320] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] ? 1'h0 : _filtered_keep_10_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[353:352] == 2'h3 & io_xbar_in_bits_tdata[353:352] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] ? 1'h0 : _filtered_keep_11_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[385:384] == 2'h3 & io_xbar_in_bits_tdata[385:384] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] ? 1'h0 : _filtered_keep_12_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[417:416] == 2'h3 & io_xbar_in_bits_tdata[417:416] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] ? 1'h0 : _filtered_keep_13_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[449:448] == 2'h3 & io_xbar_in_bits_tdata[449:448] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] ? 1'h0 : _filtered_keep_14_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[bfs_remote.scala 306:15]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[481:480] == 2'h3 & io_xbar_in_bits_tdata[481:480] != local_fpga_id
    ; // @[bfs_remote.scala 300:52]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] ? 1'h0 : _filtered_keep_15_T_8; // @[bfs_remote.scala 307:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[bfs_remote.scala 306:15]
  wire [7:0] collector_io_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[bfs_remote.scala 314:53]
  wire [7:0] collector_io_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[bfs_remote.scala 314:53]
  reg [31:0] vertex_in_fifo_data_count; // @[bfs_remote.scala 320:42]
  wire  _T_1 = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 321:90]
  wire  _T_2 = vertex_in_fifo_s_axis_tvalid & vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 321:49]
  wire  _T_3 = vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 322:44]
  wire  _T_5 = vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 322:88]
  wire [31:0] _vertex_in_fifo_data_count_T_1 = vertex_in_fifo_data_count + 32'h1; // @[bfs_remote.scala 325:60]
  wire [31:0] _vertex_in_fifo_data_count_T_3 = vertex_in_fifo_data_count - 32'h1; // @[bfs_remote.scala 327:60]
  reg [2:0] sync_status; // @[bfs_remote.scala 345:28]
  reg [31:0] stall_time; // @[bfs_remote.scala 346:27]
  wire  _T_13 = sync_status == 3'h6; // @[bfs_remote.scala 348:20]
  wire [31:0] _stall_time_T_1 = stall_time + 32'h1; // @[bfs_remote.scala 349:30]
  wire  _T_21 = sync_status == 3'h1; // @[bfs_remote.scala 357:26]
  wire  _T_29 = sync_status == 3'h3; // @[bfs_remote.scala 363:26]
  wire [2:0] _GEN_4 = sync_status == 3'h4 & io_signal ? 3'h0 : sync_status; // @[bfs_remote.scala 365:58 bfs_remote.scala 366:17 bfs_remote.scala 345:28]
  wire [2:0] _GEN_5 = sync_status == 3'h3 & _T_1 ? 3'h4 : _GEN_4; // @[bfs_remote.scala 363:95 bfs_remote.scala 364:17]
  wire [2:0] _GEN_6 = _T_13 & stall_time == 32'h1e ? 3'h3 : _GEN_5; // @[bfs_remote.scala 361:71 bfs_remote.scala 362:17]
  wire [2:0] _GEN_7 = sync_status == 3'h2 & io_recv_sync_phase2 ? 3'h6 : _GEN_6; // @[bfs_remote.scala 359:73 bfs_remote.scala 360:17]
  wire  need_to_send_sync = _T_21 | _T_29; // @[bfs_remote.scala 372:66]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = need_to_send_sync ? 16'h1 : collector_io_out_bits_tkeep; // @[bfs_remote.scala 376:40]
  wire [3:0] sync_data_level = level[3:0]; // @[bfs_remote.scala 339:23 bfs_remote.scala 342:19]
  wire [31:0] _vertex_in_fifo_io_s_axis_tdata_T = {1'h1,local_fpga_id,sync_data_level,25'h0}; // @[bfs_remote.scala 378:76]
  reg [31:0] send_count; // @[bfs_remote.scala 382:27]
  reg [31:0] pending_time; // @[bfs_remote.scala 383:29]
  reg [31:0] extra_time; // @[bfs_remote.scala 384:27]
  wire [31:0] _io_remote_out_bits_tlast_T_1 = packet_size - 32'h1; // @[bfs_remote.scala 389:59]
  wire  _io_remote_out_bits_tlast_T_2 = send_count == _io_remote_out_bits_tlast_T_1; // @[bfs_remote.scala 389:42]
  wire  _flow_control_unit_io_handshake_T = io_remote_out_valid & io_remote_out_ready; // @[bfs_remote.scala 392:57]
  wire  _T_34 = pending_time == 32'h0; // @[bfs_remote.scala 399:27]
  wire [31:0] _extra_time_T_1 = extra_time + 32'h1; // @[bfs_remote.scala 400:30]
  wire [31:0] _pending_time_T_2 = flow_control_unit_io_pending_bits - extra_time; // @[bfs_remote.scala 406:46]
  wire [31:0] _pending_time_T_5 = pending_time - 32'h1; // @[bfs_remote.scala 408:34]
  wire [31:0] _send_count_T_1 = send_count + 32'h1; // @[bfs_remote.scala 414:32]
  wire  _T_42 = vertex_in_fifo_data_count >= packet_size & send_count == 32'h0; // @[bfs_remote.scala 417:49]
  wire  _T_44 = _T_42 | send_count != 32'h0; // @[bfs_remote.scala 418:3]
  wire  _GEN_17 = _T_34 & vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 420:31 bfs_remote.scala 421:27 bfs_remote.scala 402:23]
  wire  _GEN_18 = _T_34 & io_remote_out_ready; // @[bfs_remote.scala 420:31 bfs_remote.scala 422:39 bfs_remote.scala 403:35]
  axis_data_collector collector ( // @[bfs_remote.scala 312:25]
    .clock(collector_clock),
    .reset(collector_reset),
    .io_in_ready(collector_io_in_ready),
    .io_in_valid(collector_io_in_valid),
    .io_in_bits_tdata(collector_io_in_bits_tdata),
    .io_in_bits_tkeep(collector_io_in_bits_tkeep),
    .io_out_ready(collector_io_out_ready),
    .io_out_valid(collector_io_out_valid),
    .io_out_bits_tdata(collector_io_out_bits_tdata),
    .io_out_bits_tkeep(collector_io_out_bits_tkeep),
    .io_out_bits_tlast(collector_io_out_bits_tlast),
    .io_flush(collector_io_flush),
    .io_empty(collector_io_empty)
  );
  remote_apply_vid_fifo vertex_in_fifo ( // @[bfs_remote.scala 319:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .axis_rd_data_count(vertex_in_fifo_axis_rd_data_count)
  );
  flow_control flow_control_unit ( // @[bfs_remote.scala 385:33]
    .clock(flow_control_unit_clock),
    .reset(flow_control_unit_reset),
    .io_data(flow_control_unit_io_data),
    .io_keep(flow_control_unit_io_keep),
    .io_handshake(flow_control_unit_io_handshake),
    .io_handshake_last(flow_control_unit_io_handshake_last),
    .io_period(flow_control_unit_io_period),
    .io_pending_valid(flow_control_unit_io_pending_valid),
    .io_pending_bits(flow_control_unit_io_pending_bits),
    .io_parameter(flow_control_unit_io_parameter),
    .io_idol_fpga_num(flow_control_unit_io_idol_fpga_num)
  );
  assign io_xbar_in_ready = collector_io_in_ready; // @[bfs_remote.scala 317:20]
  assign io_remote_out_valid = (_T_44 | sync_status != 3'h0) & _GEN_17; // @[bfs_remote.scala 419:33 bfs_remote.scala 402:23]
  assign io_remote_out_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 387:28]
  assign io_remote_out_bits_tkeep = vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 386:28]
  assign io_remote_out_bits_tlast = send_count == _io_remote_out_bits_tlast_T_1 | vertex_in_fifo_data_count == 32'h1; // @[bfs_remote.scala 389:66]
  assign io_signal_ack = sync_status == 3'h4; // @[bfs_remote.scala 368:32]
  assign io_end = _T_29 & _T_1; // @[bfs_remote.scala 369:50]
  assign collector_clock = clock;
  assign collector_reset = reset;
  assign collector_io_in_valid = io_xbar_in_valid; // @[bfs_remote.scala 313:25]
  assign collector_io_in_bits_tdata = io_xbar_in_bits_tdata; // @[bfs_remote.scala 315:30]
  assign collector_io_in_bits_tkeep = {collector_io_in_bits_tkeep_hi,collector_io_in_bits_tkeep_lo}; // @[bfs_remote.scala 314:53]
  assign collector_io_out_ready = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 379:26]
  assign collector_io_flush = sync_status == 3'h5; // @[bfs_remote.scala 370:37]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[bfs_remote.scala 373:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[bfs_remote.scala 374:39]
  assign vertex_in_fifo_s_axis_tdata = need_to_send_sync ? {{480'd0}, _vertex_in_fifo_io_s_axis_tdata_T} :
    collector_io_out_bits_tdata; // @[bfs_remote.scala 378:40]
  assign vertex_in_fifo_s_axis_tvalid = collector_io_out_valid | need_to_send_sync; // @[bfs_remote.scala 375:63]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T}; // @[bfs_remote.scala 376:40]
  assign vertex_in_fifo_s_axis_tlast = 1'h1; // @[bfs_remote.scala 377:34]
  assign vertex_in_fifo_m_axis_tready = (_T_44 | sync_status != 3'h0) & _GEN_18; // @[bfs_remote.scala 419:33 bfs_remote.scala 403:35]
  assign flow_control_unit_clock = clock;
  assign flow_control_unit_reset = reset;
  assign flow_control_unit_io_data = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 390:29]
  assign flow_control_unit_io_keep = vertex_in_fifo_m_axis_tkeep[15:0]; // @[bfs_remote.scala 391:29]
  assign flow_control_unit_io_handshake = io_remote_out_valid & io_remote_out_ready; // @[bfs_remote.scala 392:57]
  assign flow_control_unit_io_handshake_last = io_remote_out_bits_tlast; // @[bfs_remote.scala 393:39]
  assign flow_control_unit_io_period = pending_period; // @[bfs_remote.scala 394:31]
  assign flow_control_unit_io_parameter = pending_parameter; // @[bfs_remote.scala 395:34]
  assign flow_control_unit_io_idol_fpga_num = io_idol_fpga_num; // @[bfs_remote.scala 396:38]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 288:22]
      level <= 32'h0; // @[bfs_remote.scala 288:22]
    end else begin
      level <= io_level; // @[bfs_remote.scala 289:9]
    end
    if (reset) begin // @[bfs_remote.scala 290:30]
      local_fpga_id <= 2'h0; // @[bfs_remote.scala 290:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[bfs_remote.scala 291:17]
    end
    if (reset) begin // @[bfs_remote.scala 292:28]
      packet_size <= 32'h0; // @[bfs_remote.scala 292:28]
    end else begin
      packet_size <= io_packet_size; // @[bfs_remote.scala 293:15]
    end
    if (reset) begin // @[bfs_remote.scala 294:31]
      pending_period <= 32'h0; // @[bfs_remote.scala 294:31]
    end else begin
      pending_period <= io_pending_time; // @[bfs_remote.scala 295:18]
    end
    if (reset) begin // @[bfs_remote.scala 296:34]
      pending_parameter <= 32'h0; // @[bfs_remote.scala 296:34]
    end else begin
      pending_parameter <= io_pending_parameter; // @[bfs_remote.scala 297:21]
    end
    if (reset) begin // @[bfs_remote.scala 320:42]
      vertex_in_fifo_data_count <= 32'h0; // @[bfs_remote.scala 320:42]
    end else if (!(_T_2 & vertex_in_fifo_m_axis_tvalid & vertex_in_fifo_m_axis_tready)) begin // @[bfs_remote.scala 322:92]
      if (_T_2) begin // @[bfs_remote.scala 324:99]
        vertex_in_fifo_data_count <= _vertex_in_fifo_data_count_T_1; // @[bfs_remote.scala 325:31]
      end else if (_T_3 & _T_5) begin // @[bfs_remote.scala 326:99]
        vertex_in_fifo_data_count <= _vertex_in_fifo_data_count_T_3; // @[bfs_remote.scala 327:31]
      end
    end
    if (reset) begin // @[bfs_remote.scala 345:28]
      sync_status <= 3'h0; // @[bfs_remote.scala 345:28]
    end else if (sync_status == 3'h0 & &io_recv_sync & local_fpga_id != 2'h3) begin // @[bfs_remote.scala 353:90]
      sync_status <= 3'h5; // @[bfs_remote.scala 354:17]
    end else if (sync_status == 3'h5 & collector_io_empty) begin // @[bfs_remote.scala 355:61]
      sync_status <= 3'h1; // @[bfs_remote.scala 356:17]
    end else if (sync_status == 3'h1 & _T_1) begin // @[bfs_remote.scala 357:95]
      sync_status <= 3'h2; // @[bfs_remote.scala 358:17]
    end else begin
      sync_status <= _GEN_7;
    end
    if (reset) begin // @[bfs_remote.scala 346:27]
      stall_time <= 32'h0; // @[bfs_remote.scala 346:27]
    end else if (sync_status == 3'h6) begin // @[bfs_remote.scala 348:42]
      stall_time <= _stall_time_T_1; // @[bfs_remote.scala 349:16]
    end else begin
      stall_time <= 32'h0; // @[bfs_remote.scala 351:16]
    end
    if (reset) begin // @[bfs_remote.scala 382:27]
      send_count <= 32'h0; // @[bfs_remote.scala 382:27]
    end else if (_flow_control_unit_io_handshake_T) begin // @[bfs_remote.scala 410:51]
      if (_io_remote_out_bits_tlast_T_2) begin // @[bfs_remote.scala 411:45]
        send_count <= 32'h0; // @[bfs_remote.scala 412:18]
      end else begin
        send_count <= _send_count_T_1; // @[bfs_remote.scala 414:18]
      end
    end
    if (reset) begin // @[bfs_remote.scala 383:29]
      pending_time <= 32'h0; // @[bfs_remote.scala 383:29]
    end else if (flow_control_unit_io_pending_valid) begin // @[bfs_remote.scala 404:43]
      if (extra_time > flow_control_unit_io_pending_bits) begin // @[bfs_remote.scala 405:24]
        pending_time <= 32'h0;
      end else begin
        pending_time <= _pending_time_T_2;
      end
    end else if (pending_time != 32'h0) begin // @[bfs_remote.scala 407:35]
      pending_time <= _pending_time_T_5; // @[bfs_remote.scala 408:18]
    end
    if (reset) begin // @[bfs_remote.scala 384:27]
      extra_time <= 32'h0; // @[bfs_remote.scala 384:27]
    end else if (flow_control_unit_io_pending_valid) begin // @[bfs_remote.scala 397:43]
      extra_time <= 32'h0; // @[bfs_remote.scala 398:16]
    end else if (pending_time == 32'h0) begin // @[bfs_remote.scala 399:35]
      extra_time <= _extra_time_T_1; // @[bfs_remote.scala 400:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  level = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  local_fpga_id = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  packet_size = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  pending_period = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pending_parameter = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  vertex_in_fifo_data_count = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  sync_status = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  stall_time = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  send_count = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  pending_time = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  extra_time = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Remote_Scatter(
  input          clock,
  input          reset,
  output         io_remote_in_w_ready,
  input          io_remote_in_w_valid,
  input  [511:0] io_remote_in_w_bits_wdata,
  input  [63:0]  io_remote_in_w_bits_wstrb,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [511:0] io_xbar_out_bits_tdata,
  output [15:0]  io_xbar_out_bits_tkeep,
  input          io_signal,
  input          io_start,
  output         io_issue_sync,
  output         io_issue_sync_phase2_0,
  output         io_issue_sync_phase2_1,
  output         io_issue_sync_phase2_2,
  output         io_issue_sync_phase2_3,
  input  [1:0]   io_local_fpga_id,
  output [1:0]   io_idol_fpga_num
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_in_fifo_s_axis_aclk; // @[bfs_remote.scala 550:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[bfs_remote.scala 550:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[bfs_remote.scala 550:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[bfs_remote.scala 550:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[bfs_remote.scala 550:30]
  wire  vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 550:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 550:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 550:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 550:30]
  wire  vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 550:30]
  reg [1:0] local_fpga_id; // @[bfs_remote.scala 541:30]
  wire [1:0] sync_data_id = vertex_in_fifo_m_axis_tdata[30:29]; // @[bfs_remote.scala 558:65]
  wire  sync_data_flag = vertex_in_fifo_m_axis_tdata[31]; // @[bfs_remote.scala 558:65]
  reg [3:0] syncs_0; // @[bfs_remote.scala 559:22]
  reg [3:0] syncs_1; // @[bfs_remote.scala 559:22]
  reg [3:0] syncs_2; // @[bfs_remote.scala 559:22]
  reg [3:0] syncs_3; // @[bfs_remote.scala 559:22]
  wire  _is_sync_T_4 = vertex_in_fifo_m_axis_tvalid & sync_data_flag & vertex_in_fifo_m_axis_tkeep[0]; // @[bfs_remote.scala 560:76]
  wire  is_sync = _is_sync_T_4 & ~io_issue_sync; // @[bfs_remote.scala 561:47]
  wire [3:0] _syncs_0_T_1 = syncs_0 + 4'h1; // @[bfs_remote.scala 567:22]
  wire [3:0] _syncs_1_T_1 = syncs_1 + 4'h1; // @[bfs_remote.scala 567:22]
  wire [3:0] _syncs_2_T_1 = syncs_2 + 4'h1; // @[bfs_remote.scala 567:22]
  wire [3:0] _syncs_3_T_1 = syncs_3 + 4'h1; // @[bfs_remote.scala 567:22]
  wire  _T_32 = syncs_0 > 4'h0; // @[bfs_remote.scala 573:70]
  wire  _T_33 = syncs_1 > 4'h0; // @[bfs_remote.scala 573:70]
  wire  _T_34 = syncs_2 > 4'h0; // @[bfs_remote.scala 573:70]
  wire  _T_35 = syncs_3 > 4'h0; // @[bfs_remote.scala 573:70]
  wire [3:0] _io_idol_fpga_num_WIRE = {{3'd0}, _T_32}; // @[bfs_remote.scala 575:54 bfs_remote.scala 575:54]
  wire [3:0] _io_idol_fpga_num_WIRE_1 = {{3'd0}, _T_33}; // @[bfs_remote.scala 575:54 bfs_remote.scala 575:54]
  wire [3:0] _io_idol_fpga_num_T_5 = _io_idol_fpga_num_WIRE + _io_idol_fpga_num_WIRE_1; // @[bfs_remote.scala 575:82]
  wire [3:0] _io_idol_fpga_num_WIRE_2 = {{3'd0}, _T_34}; // @[bfs_remote.scala 575:54 bfs_remote.scala 575:54]
  wire [3:0] _io_idol_fpga_num_T_7 = _io_idol_fpga_num_T_5 + _io_idol_fpga_num_WIRE_2; // @[bfs_remote.scala 575:82]
  wire [3:0] _io_idol_fpga_num_WIRE_3 = {{3'd0}, _T_35}; // @[bfs_remote.scala 575:54 bfs_remote.scala 575:54]
  wire [3:0] _io_idol_fpga_num_T_9 = _io_idol_fpga_num_T_7 + _io_idol_fpga_num_WIRE_3; // @[bfs_remote.scala 575:82]
  wire [3:0] _io_idol_fpga_num_T_11 = _io_idol_fpga_num_T_9 - 4'h1; // @[bfs_remote.scala 575:86]
  wire [63:0] _io_xbar_out_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 143:21]
  wire  _io_xbar_out_valid_T = is_sync ? 1'h0 : vertex_in_fifo_m_axis_tvalid; // @[Mux.scala 98:16]
  reg [31:0] packet_recv; // @[bfs_remote.scala 598:28]
  wire [31:0] _packet_recv_T_1 = packet_recv + 32'h1; // @[bfs_remote.scala 601:32]
  reg [31:0] ready_counter; // @[bfs_remote.scala 604:30]
  wire [31:0] _ready_counter_T_1 = ready_counter + 32'h1; // @[bfs_remote.scala 607:36]
  remote_vid_fifo vertex_in_fifo ( // @[bfs_remote.scala 550:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready)
  );
  assign io_remote_in_w_ready = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 556:24]
  assign io_xbar_out_valid = io_issue_sync ? 1'h0 : _io_xbar_out_valid_T; // @[Mux.scala 98:16]
  assign io_xbar_out_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 142:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 143:13]
  assign io_issue_sync = syncs_0 == 4'h2 & syncs_1 == 4'h2 & syncs_2 == 4'h2 & syncs_3 == 4'h2; // @[bfs_remote.scala 574:54]
  assign io_issue_sync_phase2_0 = syncs_0 > 4'h0 & syncs_1 > 4'h0 & syncs_2 > 4'h0 & syncs_3 > 4'h0; // @[bfs_remote.scala 573:86]
  assign io_issue_sync_phase2_1 = syncs_0 > 4'h0 & syncs_1 > 4'h0 & syncs_2 > 4'h0 & syncs_3 > 4'h0; // @[bfs_remote.scala 573:86]
  assign io_issue_sync_phase2_2 = syncs_0 > 4'h0 & syncs_1 > 4'h0 & syncs_2 > 4'h0 & syncs_3 > 4'h0; // @[bfs_remote.scala 573:86]
  assign io_issue_sync_phase2_3 = syncs_0 > 4'h0 & syncs_1 > 4'h0 & syncs_2 > 4'h0 & syncs_3 > 4'h0; // @[bfs_remote.scala 573:86]
  assign io_idol_fpga_num = _io_idol_fpga_num_T_11[1:0]; // @[bfs_remote.scala 575:20]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[bfs_remote.scala 551:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[bfs_remote.scala 552:39]
  assign vertex_in_fifo_s_axis_tdata = io_remote_in_w_bits_wdata; // @[bfs_remote.scala 555:34]
  assign vertex_in_fifo_s_axis_tvalid = io_remote_in_w_valid; // @[bfs_remote.scala 553:35]
  assign vertex_in_fifo_s_axis_tkeep = io_remote_in_w_bits_wstrb; // @[bfs_remote.scala 554:34]
  assign vertex_in_fifo_m_axis_tready = io_issue_sync ? 1'h0 : is_sync | io_xbar_out_ready; // @[Mux.scala 98:16]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 541:30]
      local_fpga_id <= 2'h0; // @[bfs_remote.scala 541:30]
    end else begin
      local_fpga_id <= io_local_fpga_id; // @[bfs_remote.scala 542:17]
    end
    if (reset) begin // @[bfs_remote.scala 559:22]
      syncs_0 <= 4'h0; // @[bfs_remote.scala 559:22]
    end else if (local_fpga_id == 2'h0 & io_start) begin // @[bfs_remote.scala 564:46]
      syncs_0 <= 4'h2; // @[bfs_remote.scala 565:14]
    end else if (is_sync & sync_data_id == 2'h0) begin // @[bfs_remote.scala 566:50]
      syncs_0 <= _syncs_0_T_1; // @[bfs_remote.scala 567:14]
    end else if (~io_start & io_signal & local_fpga_id != 2'h0) begin // @[bfs_remote.scala 568:66]
      syncs_0 <= 4'h0; // @[bfs_remote.scala 569:14]
    end
    if (reset) begin // @[bfs_remote.scala 559:22]
      syncs_1 <= 4'h0; // @[bfs_remote.scala 559:22]
    end else if (local_fpga_id == 2'h1 & io_start) begin // @[bfs_remote.scala 564:46]
      syncs_1 <= 4'h2; // @[bfs_remote.scala 565:14]
    end else if (is_sync & sync_data_id == 2'h1) begin // @[bfs_remote.scala 566:50]
      syncs_1 <= _syncs_1_T_1; // @[bfs_remote.scala 567:14]
    end else if (~io_start & io_signal & local_fpga_id != 2'h1) begin // @[bfs_remote.scala 568:66]
      syncs_1 <= 4'h0; // @[bfs_remote.scala 569:14]
    end
    if (reset) begin // @[bfs_remote.scala 559:22]
      syncs_2 <= 4'h0; // @[bfs_remote.scala 559:22]
    end else if (local_fpga_id == 2'h2 & io_start) begin // @[bfs_remote.scala 564:46]
      syncs_2 <= 4'h2; // @[bfs_remote.scala 565:14]
    end else if (is_sync & sync_data_id == 2'h2) begin // @[bfs_remote.scala 566:50]
      syncs_2 <= _syncs_2_T_1; // @[bfs_remote.scala 567:14]
    end else if (~io_start & io_signal & local_fpga_id != 2'h2) begin // @[bfs_remote.scala 568:66]
      syncs_2 <= 4'h0; // @[bfs_remote.scala 569:14]
    end
    if (reset) begin // @[bfs_remote.scala 559:22]
      syncs_3 <= 4'h0; // @[bfs_remote.scala 559:22]
    end else if (local_fpga_id == 2'h3 & io_start) begin // @[bfs_remote.scala 564:46]
      syncs_3 <= 4'h2; // @[bfs_remote.scala 565:14]
    end else if (is_sync & sync_data_id == 2'h3) begin // @[bfs_remote.scala 566:50]
      syncs_3 <= _syncs_3_T_1; // @[bfs_remote.scala 567:14]
    end else if (~io_start & io_signal & local_fpga_id != 2'h3) begin // @[bfs_remote.scala 568:66]
      syncs_3 <= 4'h0; // @[bfs_remote.scala 569:14]
    end
    if (reset) begin // @[bfs_remote.scala 598:28]
      packet_recv <= 32'h0; // @[bfs_remote.scala 598:28]
    end else if (io_remote_in_w_valid & io_remote_in_w_ready) begin // @[bfs_remote.scala 600:53]
      packet_recv <= _packet_recv_T_1; // @[bfs_remote.scala 601:17]
    end
    if (reset) begin // @[bfs_remote.scala 604:30]
      ready_counter <= 32'h0; // @[bfs_remote.scala 604:30]
    end else if (io_remote_in_w_valid & ~io_remote_in_w_ready) begin // @[bfs_remote.scala 606:65]
      ready_counter <= _ready_counter_T_1; // @[bfs_remote.scala 607:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  local_fpga_id = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  syncs_0 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  syncs_1 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  syncs_2 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  syncs_3 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  packet_recv = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  ready_counter = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_to_axi(
  input          clock,
  input          reset,
  output         io_xbar_in_0_ready,
  input          io_xbar_in_0_valid,
  input  [511:0] io_xbar_in_0_bits_tdata,
  input  [63:0]  io_xbar_in_0_bits_tkeep,
  input          io_xbar_in_0_bits_tlast,
  output         io_xbar_in_1_ready,
  input          io_xbar_in_1_valid,
  input  [511:0] io_xbar_in_1_bits_tdata,
  input  [63:0]  io_xbar_in_1_bits_tkeep,
  input          io_xbar_in_1_bits_tlast,
  output         io_xbar_in_2_ready,
  input          io_xbar_in_2_valid,
  input  [511:0] io_xbar_in_2_bits_tdata,
  input  [63:0]  io_xbar_in_2_bits_tkeep,
  input          io_xbar_in_2_bits_tlast,
  output         io_xbar_in_3_ready,
  input          io_xbar_in_3_valid,
  input  [511:0] io_xbar_in_3_bits_tdata,
  input  [63:0]  io_xbar_in_3_bits_tkeep,
  input          io_xbar_in_3_bits_tlast,
  input          io_remote_out_aw_ready,
  output         io_remote_out_aw_valid,
  output [63:0]  io_remote_out_aw_bits_awaddr,
  input          io_remote_out_w_ready,
  output         io_remote_out_w_valid,
  output [511:0] io_remote_out_w_bits_wdata,
  output [63:0]  io_remote_out_w_bits_wstrb,
  output         io_remote_out_w_bits_wlast,
  input  [63:0]  io_level_base_addr_0,
  input  [63:0]  io_level_base_addr_1,
  input  [63:0]  io_level_base_addr_2,
  input  [63:0]  io_level_base_addr_3,
  input  [31:0]  io_net_constrain
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  switch_aclk; // @[bfs_remote.scala 443:22]
  wire  switch_aresetn; // @[bfs_remote.scala 443:22]
  wire [2047:0] switch_s_axis_tdata; // @[bfs_remote.scala 443:22]
  wire [3:0] switch_s_axis_tvalid; // @[bfs_remote.scala 443:22]
  wire [255:0] switch_s_axis_tkeep; // @[bfs_remote.scala 443:22]
  wire [3:0] switch_s_axis_tready; // @[bfs_remote.scala 443:22]
  wire [3:0] switch_s_axis_tlast; // @[bfs_remote.scala 443:22]
  wire [7:0] switch_s_axis_tuser; // @[bfs_remote.scala 443:22]
  wire [511:0] switch_m_axis_tdata; // @[bfs_remote.scala 443:22]
  wire  switch_m_axis_tvalid; // @[bfs_remote.scala 443:22]
  wire [63:0] switch_m_axis_tkeep; // @[bfs_remote.scala 443:22]
  wire  switch_m_axis_tready; // @[bfs_remote.scala 443:22]
  wire  switch_m_axis_tlast; // @[bfs_remote.scala 443:22]
  wire [1:0] switch_m_axis_tuser; // @[bfs_remote.scala 443:22]
  wire [3:0] switch_s_req_suppress; // @[bfs_remote.scala 443:22]
  wire  vertex_in_fifo_s_axis_aclk; // @[bfs_remote.scala 456:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[bfs_remote.scala 456:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[bfs_remote.scala 456:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[bfs_remote.scala 456:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[bfs_remote.scala 456:30]
  wire  vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 456:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[bfs_remote.scala 456:30]
  wire [1:0] vertex_in_fifo_s_axis_tuser; // @[bfs_remote.scala 456:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 456:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 456:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 456:30]
  wire  vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 456:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[bfs_remote.scala 456:30]
  wire [1:0] vertex_in_fifo_m_axis_tuser; // @[bfs_remote.scala 456:30]
  reg [31:0] net_constrain; // @[bfs_remote.scala 438:30]
  wire [1:0] switch_io_s_axis_tvalid_lo = {io_xbar_in_1_valid,io_xbar_in_0_valid}; // @[bfs_remote.scala 447:72]
  wire [1:0] switch_io_s_axis_tvalid_hi = {io_xbar_in_3_valid,io_xbar_in_2_valid}; // @[bfs_remote.scala 447:72]
  wire [1023:0] switch_io_s_axis_tdata_lo = {io_xbar_in_1_bits_tdata,io_xbar_in_0_bits_tdata}; // @[bfs_remote.scala 448:76]
  wire [1023:0] switch_io_s_axis_tdata_hi = {io_xbar_in_3_bits_tdata,io_xbar_in_2_bits_tdata}; // @[bfs_remote.scala 448:76]
  wire [127:0] switch_io_s_axis_tkeep_lo = {io_xbar_in_1_bits_tkeep,io_xbar_in_0_bits_tkeep}; // @[bfs_remote.scala 449:76]
  wire [127:0] switch_io_s_axis_tkeep_hi = {io_xbar_in_3_bits_tkeep,io_xbar_in_2_bits_tkeep}; // @[bfs_remote.scala 449:76]
  wire [1:0] switch_io_s_axis_tlast_lo = {io_xbar_in_1_bits_tlast,io_xbar_in_0_bits_tlast}; // @[bfs_remote.scala 450:76]
  wire [1:0] switch_io_s_axis_tlast_hi = {io_xbar_in_3_bits_tlast,io_xbar_in_2_bits_tlast}; // @[bfs_remote.scala 450:76]
  reg [1:0] send_status; // @[bfs_remote.scala 469:28]
  wire  addr_issue = io_remote_out_aw_valid & io_remote_out_aw_ready; // @[bfs_remote.scala 470:43]
  wire  data_issue = io_remote_out_w_valid & io_remote_out_w_ready & io_remote_out_w_bits_wlast; // @[bfs_remote.scala 471:67]
  reg [31:0] BW_net_constrain; // @[bfs_remote.scala 472:33]
  wire  ready_to_issue = send_status == 2'h0 & vertex_in_fifo_m_axis_tvalid & BW_net_constrain == 32'h0; // @[bfs_remote.scala 473:93]
  wire [31:0] _BW_net_constrain_T_1 = net_constrain - 32'h1; // @[bfs_remote.scala 475:39]
  wire [31:0] _BW_net_constrain_T_3 = BW_net_constrain - 32'h1; // @[bfs_remote.scala 477:42]
  wire  _T_1 = send_status == 2'h1; // @[bfs_remote.scala 481:27]
  wire  _T_2 = send_status == 2'h1 & addr_issue; // @[bfs_remote.scala 481:42]
  wire  _T_3 = send_status == 2'h1 & addr_issue & data_issue; // @[bfs_remote.scala 481:56]
  wire  _T_4 = send_status == 2'h2; // @[bfs_remote.scala 482:21]
  wire  _T_5 = send_status == 2'h2 & addr_issue; // @[bfs_remote.scala 482:36]
  wire  _T_6 = _T_3 | send_status == 2'h2 & addr_issue; // @[bfs_remote.scala 482:5]
  wire  _T_7 = send_status == 2'h3; // @[bfs_remote.scala 483:21]
  wire [1:0] _GEN_2 = _T_2 & ~data_issue ? 2'h3 : send_status; // @[bfs_remote.scala 487:70 bfs_remote.scala 488:17 bfs_remote.scala 469:28]
  wire  _io_remote_out_aw_bits_awaddr_T = vertex_in_fifo_m_axis_tuser == 2'h0; // @[bfs_remote.scala 510:42]
  wire  _io_remote_out_aw_bits_awaddr_T_1 = vertex_in_fifo_m_axis_tuser == 2'h1; // @[bfs_remote.scala 510:42]
  wire  _io_remote_out_aw_bits_awaddr_T_2 = vertex_in_fifo_m_axis_tuser == 2'h2; // @[bfs_remote.scala 510:42]
  wire  _io_remote_out_aw_bits_awaddr_T_3 = vertex_in_fifo_m_axis_tuser == 2'h3; // @[bfs_remote.scala 510:42]
  wire [63:0] _io_remote_out_aw_bits_awaddr_T_4 = _io_remote_out_aw_bits_awaddr_T ? io_level_base_addr_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _io_remote_out_aw_bits_awaddr_T_5 = _io_remote_out_aw_bits_awaddr_T_1 ? io_level_base_addr_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _io_remote_out_aw_bits_awaddr_T_6 = _io_remote_out_aw_bits_awaddr_T_2 ? io_level_base_addr_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _io_remote_out_aw_bits_awaddr_T_7 = _io_remote_out_aw_bits_awaddr_T_3 ? io_level_base_addr_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _io_remote_out_aw_bits_awaddr_T_8 = _io_remote_out_aw_bits_awaddr_T_4 | _io_remote_out_aw_bits_awaddr_T_5; // @[Mux.scala 27:72]
  wire [63:0] _io_remote_out_aw_bits_awaddr_T_9 = _io_remote_out_aw_bits_awaddr_T_8 | _io_remote_out_aw_bits_awaddr_T_6; // @[Mux.scala 27:72]
  reg [31:0] packet_sent; // @[bfs_remote.scala 518:28]
  wire [31:0] _packet_sent_T_1 = packet_sent + 32'h1; // @[bfs_remote.scala 521:32]
  axis_to_axi_switch switch ( // @[bfs_remote.scala 443:22]
    .aclk(switch_aclk),
    .aresetn(switch_aresetn),
    .s_axis_tdata(switch_s_axis_tdata),
    .s_axis_tvalid(switch_s_axis_tvalid),
    .s_axis_tkeep(switch_s_axis_tkeep),
    .s_axis_tready(switch_s_axis_tready),
    .s_axis_tlast(switch_s_axis_tlast),
    .s_axis_tuser(switch_s_axis_tuser),
    .m_axis_tdata(switch_m_axis_tdata),
    .m_axis_tvalid(switch_m_axis_tvalid),
    .m_axis_tkeep(switch_m_axis_tkeep),
    .m_axis_tready(switch_m_axis_tready),
    .m_axis_tlast(switch_m_axis_tlast),
    .m_axis_tuser(switch_m_axis_tuser),
    .s_req_suppress(switch_s_req_suppress)
  );
  remote_vid_user_fifo vertex_in_fifo ( // @[bfs_remote.scala 456:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tuser(vertex_in_fifo_s_axis_tuser),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tuser(vertex_in_fifo_m_axis_tuser)
  );
  assign io_xbar_in_0_ready = switch_s_axis_tready[0]; // @[bfs_remote.scala 453:56]
  assign io_xbar_in_1_ready = switch_s_axis_tready[1]; // @[bfs_remote.scala 453:56]
  assign io_xbar_in_2_ready = switch_s_axis_tready[2]; // @[bfs_remote.scala 453:56]
  assign io_xbar_in_3_ready = switch_s_axis_tready[3]; // @[bfs_remote.scala 453:56]
  assign io_remote_out_aw_valid = _T_1 | _T_4; // @[bfs_remote.scala 503:56]
  assign io_remote_out_aw_bits_awaddr = _io_remote_out_aw_bits_awaddr_T_9 | _io_remote_out_aw_bits_awaddr_T_7; // @[Mux.scala 27:72]
  assign io_remote_out_w_valid = _T_1 | _T_7; // @[bfs_remote.scala 513:55]
  assign io_remote_out_w_bits_wdata = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 515:30]
  assign io_remote_out_w_bits_wstrb = {{48'd0}, vertex_in_fifo_m_axis_tkeep[15:0]}; // @[bfs_remote.scala 516:63]
  assign io_remote_out_w_bits_wlast = vertex_in_fifo_m_axis_tlast; // @[bfs_remote.scala 514:30]
  assign switch_aclk = clock; // @[bfs_remote.scala 444:33]
  assign switch_aresetn = ~reset; // @[bfs_remote.scala 445:24]
  assign switch_s_axis_tdata = {switch_io_s_axis_tdata_hi,switch_io_s_axis_tdata_lo}; // @[bfs_remote.scala 448:76]
  assign switch_s_axis_tvalid = {switch_io_s_axis_tvalid_hi,switch_io_s_axis_tvalid_lo}; // @[bfs_remote.scala 447:72]
  assign switch_s_axis_tkeep = {switch_io_s_axis_tkeep_hi,switch_io_s_axis_tkeep_lo}; // @[bfs_remote.scala 449:76]
  assign switch_s_axis_tlast = {switch_io_s_axis_tlast_hi,switch_io_s_axis_tlast_lo}; // @[bfs_remote.scala 450:76]
  assign switch_s_axis_tuser = 8'he4; // @[bfs_remote.scala 451:76]
  assign switch_m_axis_tready = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 460:28]
  assign switch_s_req_suppress = 4'h0; // @[bfs_remote.scala 446:28]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[bfs_remote.scala 458:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[bfs_remote.scala 459:39]
  assign vertex_in_fifo_s_axis_tdata = switch_m_axis_tdata; // @[bfs_remote.scala 460:28]
  assign vertex_in_fifo_s_axis_tvalid = switch_m_axis_tvalid; // @[bfs_remote.scala 460:28]
  assign vertex_in_fifo_s_axis_tkeep = switch_m_axis_tkeep; // @[bfs_remote.scala 460:28]
  assign vertex_in_fifo_s_axis_tlast = switch_m_axis_tlast; // @[bfs_remote.scala 460:28]
  assign vertex_in_fifo_s_axis_tuser = switch_m_axis_tuser; // @[bfs_remote.scala 460:28]
  assign vertex_in_fifo_m_axis_tready = _T_1 | _T_7 ? io_remote_out_w_ready : _T_5; // @[bfs_remote.scala 491:64 bfs_remote.scala 492:37]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 438:30]
      net_constrain <= 32'h0; // @[bfs_remote.scala 438:30]
    end else begin
      net_constrain <= io_net_constrain; // @[bfs_remote.scala 439:17]
    end
    if (reset) begin // @[bfs_remote.scala 469:28]
      send_status <= 2'h0; // @[bfs_remote.scala 469:28]
    end else if (ready_to_issue) begin // @[bfs_remote.scala 479:23]
      send_status <= 2'h1; // @[bfs_remote.scala 480:17]
    end else if (_T_6 | send_status == 2'h3 & data_issue) begin // @[bfs_remote.scala 483:50]
      send_status <= 2'h0; // @[bfs_remote.scala 484:17]
    end else if (_T_1 & ~addr_issue & data_issue) begin // @[bfs_remote.scala 485:70]
      send_status <= 2'h2; // @[bfs_remote.scala 486:17]
    end else begin
      send_status <= _GEN_2;
    end
    if (reset) begin // @[bfs_remote.scala 472:33]
      BW_net_constrain <= 32'h0; // @[bfs_remote.scala 472:33]
    end else if (ready_to_issue) begin // @[bfs_remote.scala 474:23]
      BW_net_constrain <= _BW_net_constrain_T_1; // @[bfs_remote.scala 475:22]
    end else if (BW_net_constrain != 32'h0) begin // @[bfs_remote.scala 476:39]
      BW_net_constrain <= _BW_net_constrain_T_3; // @[bfs_remote.scala 477:22]
    end
    if (reset) begin // @[bfs_remote.scala 518:28]
      packet_sent <= 32'h0; // @[bfs_remote.scala 518:28]
    end else if (addr_issue) begin // @[bfs_remote.scala 520:57]
      packet_sent <= _packet_sent_T_1; // @[bfs_remote.scala 521:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  net_constrain = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  send_status = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  BW_net_constrain = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  packet_sent = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BFS_ps(
  input          clock,
  input          reset,
  input  [63:0]  io_config_awaddr,
  input          io_config_awvalid,
  output         io_config_awready,
  input  [63:0]  io_config_araddr,
  input          io_config_arvalid,
  output         io_config_arready,
  input  [31:0]  io_config_wdata,
  input  [3:0]   io_config_wstrb,
  input          io_config_wvalid,
  output         io_config_wready,
  output [31:0]  io_config_rdata,
  output [1:0]   io_config_rresp,
  output         io_config_rvalid,
  input          io_config_rready,
  output [1:0]   io_config_bresp,
  output         io_config_bvalid,
  input          io_config_bready,
  input          io_PLmemory_0_aw_ready,
  output         io_PLmemory_0_aw_valid,
  output [63:0]  io_PLmemory_0_aw_bits_awaddr,
  output [6:0]   io_PLmemory_0_aw_bits_awid,
  output [7:0]   io_PLmemory_0_aw_bits_awlen,
  output [2:0]   io_PLmemory_0_aw_bits_awsize,
  output [1:0]   io_PLmemory_0_aw_bits_awburst,
  output         io_PLmemory_0_aw_bits_awlock,
  input          io_PLmemory_0_ar_ready,
  output         io_PLmemory_0_ar_valid,
  output [63:0]  io_PLmemory_0_ar_bits_araddr,
  output [6:0]   io_PLmemory_0_ar_bits_arid,
  output [7:0]   io_PLmemory_0_ar_bits_arlen,
  output [2:0]   io_PLmemory_0_ar_bits_arsize,
  output [1:0]   io_PLmemory_0_ar_bits_arburst,
  output         io_PLmemory_0_ar_bits_arlock,
  input          io_PLmemory_0_w_ready,
  output         io_PLmemory_0_w_valid,
  output [511:0] io_PLmemory_0_w_bits_wdata,
  output [63:0]  io_PLmemory_0_w_bits_wstrb,
  output         io_PLmemory_0_w_bits_wlast,
  output         io_PLmemory_0_r_ready,
  input          io_PLmemory_0_r_valid,
  input  [511:0] io_PLmemory_0_r_bits_rdata,
  input  [6:0]   io_PLmemory_0_r_bits_rid,
  input          io_PLmemory_0_r_bits_rlast,
  output         io_PLmemory_0_b_ready,
  input          io_PLmemory_0_b_valid,
  input  [1:0]   io_PLmemory_0_b_bits_bresp,
  input  [6:0]   io_PLmemory_0_b_bits_bid,
  input          io_PLmemory_1_aw_ready,
  output         io_PLmemory_1_aw_valid,
  output [63:0]  io_PLmemory_1_aw_bits_awaddr,
  output [6:0]   io_PLmemory_1_aw_bits_awid,
  output [7:0]   io_PLmemory_1_aw_bits_awlen,
  output [2:0]   io_PLmemory_1_aw_bits_awsize,
  output [1:0]   io_PLmemory_1_aw_bits_awburst,
  output         io_PLmemory_1_aw_bits_awlock,
  input          io_PLmemory_1_ar_ready,
  output         io_PLmemory_1_ar_valid,
  output [63:0]  io_PLmemory_1_ar_bits_araddr,
  output [6:0]   io_PLmemory_1_ar_bits_arid,
  output [7:0]   io_PLmemory_1_ar_bits_arlen,
  output [2:0]   io_PLmemory_1_ar_bits_arsize,
  output [1:0]   io_PLmemory_1_ar_bits_arburst,
  output         io_PLmemory_1_ar_bits_arlock,
  input          io_PLmemory_1_w_ready,
  output         io_PLmemory_1_w_valid,
  output [511:0] io_PLmemory_1_w_bits_wdata,
  output [63:0]  io_PLmemory_1_w_bits_wstrb,
  output         io_PLmemory_1_w_bits_wlast,
  output         io_PLmemory_1_r_ready,
  input          io_PLmemory_1_r_valid,
  input  [511:0] io_PLmemory_1_r_bits_rdata,
  input  [6:0]   io_PLmemory_1_r_bits_rid,
  input          io_PLmemory_1_r_bits_rlast,
  output         io_PLmemory_1_b_ready,
  input          io_PLmemory_1_b_valid,
  input  [1:0]   io_PLmemory_1_b_bits_bresp,
  input  [6:0]   io_PLmemory_1_b_bits_bid,
  input          io_PSmemory_0_aw_ready,
  output         io_PSmemory_0_aw_valid,
  output [63:0]  io_PSmemory_0_aw_bits_awaddr,
  output [5:0]   io_PSmemory_0_aw_bits_awid,
  output [7:0]   io_PSmemory_0_aw_bits_awlen,
  output [2:0]   io_PSmemory_0_aw_bits_awsize,
  output [1:0]   io_PSmemory_0_aw_bits_awburst,
  output         io_PSmemory_0_aw_bits_awlock,
  input          io_PSmemory_0_ar_ready,
  output         io_PSmemory_0_ar_valid,
  output [63:0]  io_PSmemory_0_ar_bits_araddr,
  output [5:0]   io_PSmemory_0_ar_bits_arid,
  output [7:0]   io_PSmemory_0_ar_bits_arlen,
  output [2:0]   io_PSmemory_0_ar_bits_arsize,
  output [1:0]   io_PSmemory_0_ar_bits_arburst,
  output         io_PSmemory_0_ar_bits_arlock,
  input          io_PSmemory_0_w_ready,
  output         io_PSmemory_0_w_valid,
  output [127:0] io_PSmemory_0_w_bits_wdata,
  output [15:0]  io_PSmemory_0_w_bits_wstrb,
  output         io_PSmemory_0_w_bits_wlast,
  output         io_PSmemory_0_r_ready,
  input          io_PSmemory_0_r_valid,
  input  [127:0] io_PSmemory_0_r_bits_rdata,
  input  [5:0]   io_PSmemory_0_r_bits_rid,
  input          io_PSmemory_0_r_bits_rlast,
  output         io_PSmemory_0_b_ready,
  input          io_PSmemory_0_b_valid,
  input  [1:0]   io_PSmemory_0_b_bits_bresp,
  input  [5:0]   io_PSmemory_0_b_bits_bid,
  input          io_PSmemory_1_aw_ready,
  output         io_PSmemory_1_aw_valid,
  output [63:0]  io_PSmemory_1_aw_bits_awaddr,
  output [5:0]   io_PSmemory_1_aw_bits_awid,
  output [7:0]   io_PSmemory_1_aw_bits_awlen,
  output [2:0]   io_PSmemory_1_aw_bits_awsize,
  output [1:0]   io_PSmemory_1_aw_bits_awburst,
  output         io_PSmemory_1_aw_bits_awlock,
  input          io_PSmemory_1_ar_ready,
  output         io_PSmemory_1_ar_valid,
  output [63:0]  io_PSmemory_1_ar_bits_araddr,
  output [5:0]   io_PSmemory_1_ar_bits_arid,
  output [7:0]   io_PSmemory_1_ar_bits_arlen,
  output [2:0]   io_PSmemory_1_ar_bits_arsize,
  output [1:0]   io_PSmemory_1_ar_bits_arburst,
  output         io_PSmemory_1_ar_bits_arlock,
  input          io_PSmemory_1_w_ready,
  output         io_PSmemory_1_w_valid,
  output [127:0] io_PSmemory_1_w_bits_wdata,
  output [15:0]  io_PSmemory_1_w_bits_wstrb,
  output         io_PSmemory_1_w_bits_wlast,
  output         io_PSmemory_1_r_ready,
  input          io_PSmemory_1_r_valid,
  input  [127:0] io_PSmemory_1_r_bits_rdata,
  input  [5:0]   io_PSmemory_1_r_bits_rid,
  input          io_PSmemory_1_r_bits_rlast,
  output         io_PSmemory_1_b_ready,
  input          io_PSmemory_1_b_valid,
  input  [1:0]   io_PSmemory_1_b_bits_bresp,
  input  [5:0]   io_PSmemory_1_b_bits_bid,
  input          io_PSmemory_2_aw_ready,
  output         io_PSmemory_2_aw_valid,
  output [63:0]  io_PSmemory_2_aw_bits_awaddr,
  output [5:0]   io_PSmemory_2_aw_bits_awid,
  output [7:0]   io_PSmemory_2_aw_bits_awlen,
  output [2:0]   io_PSmemory_2_aw_bits_awsize,
  output [1:0]   io_PSmemory_2_aw_bits_awburst,
  output         io_PSmemory_2_aw_bits_awlock,
  input          io_PSmemory_2_ar_ready,
  output         io_PSmemory_2_ar_valid,
  output [63:0]  io_PSmemory_2_ar_bits_araddr,
  output [5:0]   io_PSmemory_2_ar_bits_arid,
  output [7:0]   io_PSmemory_2_ar_bits_arlen,
  output [2:0]   io_PSmemory_2_ar_bits_arsize,
  output [1:0]   io_PSmemory_2_ar_bits_arburst,
  output         io_PSmemory_2_ar_bits_arlock,
  input          io_PSmemory_2_w_ready,
  output         io_PSmemory_2_w_valid,
  output [127:0] io_PSmemory_2_w_bits_wdata,
  output [15:0]  io_PSmemory_2_w_bits_wstrb,
  output         io_PSmemory_2_w_bits_wlast,
  output         io_PSmemory_2_r_ready,
  input          io_PSmemory_2_r_valid,
  input  [127:0] io_PSmemory_2_r_bits_rdata,
  input  [5:0]   io_PSmemory_2_r_bits_rid,
  input          io_PSmemory_2_r_bits_rlast,
  output         io_PSmemory_2_b_ready,
  input          io_PSmemory_2_b_valid,
  input  [1:0]   io_PSmemory_2_b_bits_bresp,
  input  [5:0]   io_PSmemory_2_b_bits_bid,
  input          io_PSmemory_3_aw_ready,
  output         io_PSmemory_3_aw_valid,
  output [63:0]  io_PSmemory_3_aw_bits_awaddr,
  output [5:0]   io_PSmemory_3_aw_bits_awid,
  output [7:0]   io_PSmemory_3_aw_bits_awlen,
  output [2:0]   io_PSmemory_3_aw_bits_awsize,
  output [1:0]   io_PSmemory_3_aw_bits_awburst,
  output         io_PSmemory_3_aw_bits_awlock,
  input          io_PSmemory_3_ar_ready,
  output         io_PSmemory_3_ar_valid,
  output [63:0]  io_PSmemory_3_ar_bits_araddr,
  output [5:0]   io_PSmemory_3_ar_bits_arid,
  output [7:0]   io_PSmemory_3_ar_bits_arlen,
  output [2:0]   io_PSmemory_3_ar_bits_arsize,
  output [1:0]   io_PSmemory_3_ar_bits_arburst,
  output         io_PSmemory_3_ar_bits_arlock,
  input          io_PSmemory_3_w_ready,
  output         io_PSmemory_3_w_valid,
  output [127:0] io_PSmemory_3_w_bits_wdata,
  output [15:0]  io_PSmemory_3_w_bits_wstrb,
  output         io_PSmemory_3_w_bits_wlast,
  output         io_PSmemory_3_r_ready,
  input          io_PSmemory_3_r_valid,
  input  [127:0] io_PSmemory_3_r_bits_rdata,
  input  [5:0]   io_PSmemory_3_r_bits_rid,
  input          io_PSmemory_3_r_bits_rlast,
  output         io_PSmemory_3_b_ready,
  input          io_PSmemory_3_b_valid,
  input  [1:0]   io_PSmemory_3_b_bits_bresp,
  input  [5:0]   io_PSmemory_3_b_bits_bid,
  input          io_Re_memory_out_aw_ready,
  output         io_Re_memory_out_aw_valid,
  output [63:0]  io_Re_memory_out_aw_bits_awaddr,
  output [5:0]   io_Re_memory_out_aw_bits_awid,
  output [7:0]   io_Re_memory_out_aw_bits_awlen,
  output [2:0]   io_Re_memory_out_aw_bits_awsize,
  output [1:0]   io_Re_memory_out_aw_bits_awburst,
  output         io_Re_memory_out_aw_bits_awlock,
  input          io_Re_memory_out_ar_ready,
  output         io_Re_memory_out_ar_valid,
  output [63:0]  io_Re_memory_out_ar_bits_araddr,
  output [5:0]   io_Re_memory_out_ar_bits_arid,
  output [7:0]   io_Re_memory_out_ar_bits_arlen,
  output [2:0]   io_Re_memory_out_ar_bits_arsize,
  output [1:0]   io_Re_memory_out_ar_bits_arburst,
  output         io_Re_memory_out_ar_bits_arlock,
  input          io_Re_memory_out_w_ready,
  output         io_Re_memory_out_w_valid,
  output [511:0] io_Re_memory_out_w_bits_wdata,
  output [63:0]  io_Re_memory_out_w_bits_wstrb,
  output         io_Re_memory_out_w_bits_wlast,
  output         io_Re_memory_out_r_ready,
  input          io_Re_memory_out_r_valid,
  input  [511:0] io_Re_memory_out_r_bits_rdata,
  input  [5:0]   io_Re_memory_out_r_bits_rid,
  input          io_Re_memory_out_r_bits_rlast,
  output         io_Re_memory_out_b_ready,
  input          io_Re_memory_out_b_valid,
  input  [1:0]   io_Re_memory_out_b_bits_bresp,
  input  [5:0]   io_Re_memory_out_b_bits_bid,
  output         io_Re_memory_in_aw_ready,
  input          io_Re_memory_in_aw_valid,
  input  [63:0]  io_Re_memory_in_aw_bits_awaddr,
  input  [9:0]   io_Re_memory_in_aw_bits_awid,
  input  [7:0]   io_Re_memory_in_aw_bits_awlen,
  input  [2:0]   io_Re_memory_in_aw_bits_awsize,
  input  [1:0]   io_Re_memory_in_aw_bits_awburst,
  input          io_Re_memory_in_aw_bits_awlock,
  output         io_Re_memory_in_ar_ready,
  input          io_Re_memory_in_ar_valid,
  input  [63:0]  io_Re_memory_in_ar_bits_araddr,
  input  [9:0]   io_Re_memory_in_ar_bits_arid,
  input  [7:0]   io_Re_memory_in_ar_bits_arlen,
  input  [2:0]   io_Re_memory_in_ar_bits_arsize,
  input  [1:0]   io_Re_memory_in_ar_bits_arburst,
  input          io_Re_memory_in_ar_bits_arlock,
  output         io_Re_memory_in_w_ready,
  input          io_Re_memory_in_w_valid,
  input  [511:0] io_Re_memory_in_w_bits_wdata,
  input  [63:0]  io_Re_memory_in_w_bits_wstrb,
  input          io_Re_memory_in_w_bits_wlast,
  input          io_Re_memory_in_r_ready,
  output         io_Re_memory_in_r_valid,
  output [511:0] io_Re_memory_in_r_bits_rdata,
  output [9:0]   io_Re_memory_in_r_bits_rid,
  output         io_Re_memory_in_r_bits_rlast,
  input          io_Re_memory_in_b_ready,
  output         io_Re_memory_in_b_valid,
  output [1:0]   io_Re_memory_in_b_bits_bresp,
  output [9:0]   io_Re_memory_in_b_bits_bid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  controls_clock; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_reset; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_0; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_1; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_2; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_3; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_4; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_7; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_16; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_17; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_18; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_19; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_20; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_21; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_22; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_23; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_24; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_25; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_26; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_27; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_28; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_data_29; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_0; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_1; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_2; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_3; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_4; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_5; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_6; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_7; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_8; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_9; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_10; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_11; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_12; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_13; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_14; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_15; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_16; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_17; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_18; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_fin_19; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_signal; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_start; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_level; // @[nf_arm_doce_top_main.scala 30:24]
  wire [63:0] controls_io_traveled_edges; // @[nf_arm_doce_top_main.scala 30:24]
  wire [63:0] controls_io_config_awaddr; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_awvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_awready; // @[nf_arm_doce_top_main.scala 30:24]
  wire [63:0] controls_io_config_araddr; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_arvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_arready; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_config_wdata; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_wvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_wready; // @[nf_arm_doce_top_main.scala 30:24]
  wire [31:0] controls_io_config_rdata; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_rvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_rready; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_bvalid; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_config_bready; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_flush_cache; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_flush_cache_end; // @[nf_arm_doce_top_main.scala 30:24]
  wire  controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 30:24]
  wire  MemController_clock; // @[nf_arm_doce_top_main.scala 39:29]
  wire  MemController_reset; // @[nf_arm_doce_top_main.scala 39:29]
  wire  MemController_io_cacheable_out_ready; // @[nf_arm_doce_top_main.scala 39:29]
  wire  MemController_io_cacheable_out_valid; // @[nf_arm_doce_top_main.scala 39:29]
  wire [511:0] MemController_io_cacheable_out_bits_tdata; // @[nf_arm_doce_top_main.scala 39:29]
  wire [15:0] MemController_io_cacheable_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 39:29]
  wire [31:0] MemController_io_graph_scale; // @[nf_arm_doce_top_main.scala 39:29]
  wire  MemController_io_start; // @[nf_arm_doce_top_main.scala 39:29]
  wire  MemController_io_signal; // @[nf_arm_doce_top_main.scala 39:29]
  wire  MemController_io_end; // @[nf_arm_doce_top_main.scala 39:29]
  wire  MemController_io_signal_ack; // @[nf_arm_doce_top_main.scala 39:29]
  wire  Applys_0_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_0_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_0_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_0_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_0_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_0_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_0_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_0_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_0_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_1_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_1_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_1_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_1_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_1_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_1_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_1_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_1_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_1_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_2_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_2_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_2_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_2_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_2_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_2_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_2_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_2_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_2_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_3_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_3_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_3_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_3_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_3_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_3_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_3_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_3_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_3_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_4_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_4_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_4_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_4_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_4_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_4_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_4_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_4_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_4_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_4_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_5_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_5_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_5_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_5_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_5_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_5_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_5_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_5_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_5_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_5_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_6_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_6_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_6_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_6_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_6_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_6_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_6_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_6_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_6_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_6_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_7_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_7_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_7_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_7_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_7_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_7_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_7_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_7_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_7_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_7_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_8_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_8_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_8_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_8_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_8_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_8_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_8_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_8_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_8_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_8_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_9_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_9_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_9_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_9_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_9_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_9_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_9_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_9_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_9_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_9_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_10_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_10_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_10_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_10_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_10_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_10_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_10_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_10_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_10_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_10_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_11_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_11_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_11_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_11_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_11_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_11_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_11_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_11_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_11_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_11_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_12_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_12_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_12_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_12_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_12_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_12_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_12_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_12_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_12_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_12_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_13_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_13_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_13_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_13_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_13_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_13_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_13_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_13_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_13_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_13_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_14_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_14_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_14_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_14_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_14_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_14_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_14_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_14_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_14_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_14_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_15_clock; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_15_reset; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_15_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_15_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 42:16]
  wire [511:0] Applys_15_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:16]
  wire [15:0] Applys_15_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_15_io_xbar_in_bits_tlast; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Applys_15_io_end; // @[nf_arm_doce_top_main.scala 42:16]
  wire [2:0] Applys_15_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 42:16]
  wire [31:0] Applys_15_io_graph_scale; // @[nf_arm_doce_top_main.scala 42:16]
  wire  Gathers_clock; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_reset; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_ddr_in_ready; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_ddr_in_valid; // @[nf_arm_doce_top_main.scala 44:23]
  wire [511:0] Gathers_io_ddr_in_bits_tdata; // @[nf_arm_doce_top_main.scala 44:23]
  wire [15:0] Gathers_io_ddr_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_gather_out_0_ready; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_gather_out_0_valid; // @[nf_arm_doce_top_main.scala 44:23]
  wire [31:0] Gathers_io_gather_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_gather_out_1_ready; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_gather_out_1_valid; // @[nf_arm_doce_top_main.scala 44:23]
  wire [31:0] Gathers_io_gather_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_gather_out_2_ready; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_gather_out_2_valid; // @[nf_arm_doce_top_main.scala 44:23]
  wire [31:0] Gathers_io_gather_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_gather_out_3_ready; // @[nf_arm_doce_top_main.scala 44:23]
  wire  Gathers_io_gather_out_3_valid; // @[nf_arm_doce_top_main.scala 44:23]
  wire [31:0] Gathers_io_gather_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 44:23]
  wire  LevelCache_io_end; // @[nf_arm_doce_top_main.scala 45:26]
  wire  LevelCache_io_flush; // @[nf_arm_doce_top_main.scala 45:26]
  wire  Scatters_0_clock; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_reset; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_0_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 47:16]
  wire [5:0] Scatters_0_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [7:0] Scatters_0_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 47:16]
  wire [2:0] Scatters_0_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [127:0] Scatters_0_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire [5:0] Scatters_0_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [31:0] Scatters_0_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [127:0] Scatters_0_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire [3:0] Scatters_0_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_0_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_0_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_signal; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_0_io_traveled_edges; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_start; // @[nf_arm_doce_top_main.scala 47:16]
  wire [31:0] Scatters_0_io_root; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_0_io_issue_sync; // @[nf_arm_doce_top_main.scala 47:16]
  wire [4:0] Scatters_0_io_recv_sync; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_clock; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_reset; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_1_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 47:16]
  wire [5:0] Scatters_1_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [7:0] Scatters_1_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 47:16]
  wire [2:0] Scatters_1_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [127:0] Scatters_1_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire [5:0] Scatters_1_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [31:0] Scatters_1_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [127:0] Scatters_1_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire [3:0] Scatters_1_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_1_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_1_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_signal; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_1_io_traveled_edges; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_1_io_issue_sync; // @[nf_arm_doce_top_main.scala 47:16]
  wire [4:0] Scatters_1_io_recv_sync; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_clock; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_reset; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_2_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 47:16]
  wire [5:0] Scatters_2_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [7:0] Scatters_2_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 47:16]
  wire [2:0] Scatters_2_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [127:0] Scatters_2_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire [5:0] Scatters_2_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [31:0] Scatters_2_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [127:0] Scatters_2_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire [3:0] Scatters_2_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_2_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_2_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_signal; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_2_io_traveled_edges; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_2_io_issue_sync; // @[nf_arm_doce_top_main.scala 47:16]
  wire [4:0] Scatters_2_io_recv_sync; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_clock; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_reset; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_3_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 47:16]
  wire [5:0] Scatters_3_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [7:0] Scatters_3_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 47:16]
  wire [2:0] Scatters_3_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [127:0] Scatters_3_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire [5:0] Scatters_3_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [31:0] Scatters_3_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 47:16]
  wire [127:0] Scatters_3_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 47:16]
  wire [3:0] Scatters_3_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_3_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_3_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_signal; // @[nf_arm_doce_top_main.scala 47:16]
  wire [63:0] Scatters_3_io_traveled_edges; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Scatters_3_io_issue_sync; // @[nf_arm_doce_top_main.scala 47:16]
  wire [4:0] Scatters_3_io_recv_sync; // @[nf_arm_doce_top_main.scala 47:16]
  wire  Broadcaster_clock; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_reset; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_0_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_0_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [127:0] Broadcaster_io_ddr_in_0_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [3:0] Broadcaster_io_ddr_in_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_0_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_1_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_1_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [127:0] Broadcaster_io_ddr_in_1_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [3:0] Broadcaster_io_ddr_in_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_1_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_2_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_2_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [127:0] Broadcaster_io_ddr_in_2_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [3:0] Broadcaster_io_ddr_in_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_2_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_3_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_3_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [127:0] Broadcaster_io_ddr_in_3_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [3:0] Broadcaster_io_ddr_in_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_ddr_in_3_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_0_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_0_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_0_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_1_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_1_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_1_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_2_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_2_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_2_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_3_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_3_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_3_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_4_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_4_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_4_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_4_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_5_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_5_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_5_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_5_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_5_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_6_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_6_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_6_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_6_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_6_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_7_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_7_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_7_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_7_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_7_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_8_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_8_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_8_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_8_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_8_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_9_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_9_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_9_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_9_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_9_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_10_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_10_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_10_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_10_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_10_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_11_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_11_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_11_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_11_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_11_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_12_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_12_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_12_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_12_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_12_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_13_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_13_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_13_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_13_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_13_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_14_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_14_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_14_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_14_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_14_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_15_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_15_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_pe_out_15_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_pe_out_15_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_pe_out_15_bits_tlast; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_out_0_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_out_0_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_remote_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_remote_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_out_1_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_out_1_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_remote_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_remote_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_out_2_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_out_2_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_remote_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_remote_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_out_3_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_out_3_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_remote_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_remote_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_in_ready; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_remote_in_valid; // @[nf_arm_doce_top_main.scala 50:27]
  wire [511:0] Broadcaster_io_remote_in_bits_tdata; // @[nf_arm_doce_top_main.scala 50:27]
  wire [15:0] Broadcaster_io_remote_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 50:27]
  wire [1:0] Broadcaster_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_flush; // @[nf_arm_doce_top_main.scala 50:27]
  wire  Broadcaster_io_signal; // @[nf_arm_doce_top_main.scala 50:27]
  wire  ReApplys_0_clock; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_reset; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 52:16]
  wire [511:0] ReApplys_0_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 52:16]
  wire [15:0] ReApplys_0_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_io_remote_out_ready; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 52:16]
  wire [511:0] ReApplys_0_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 52:16]
  wire [63:0] ReApplys_0_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_io_remote_out_bits_tlast; // @[nf_arm_doce_top_main.scala 52:16]
  wire [3:0] ReApplys_0_io_recv_sync; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_io_recv_sync_phase2; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_io_signal; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_io_signal_ack; // @[nf_arm_doce_top_main.scala 52:16]
  wire [1:0] ReApplys_0_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_0_io_end; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_0_io_packet_size; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_0_io_level; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_0_io_pending_time; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_0_io_pending_parameter; // @[nf_arm_doce_top_main.scala 52:16]
  wire [1:0] ReApplys_0_io_idol_fpga_num; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_clock; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_reset; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 52:16]
  wire [511:0] ReApplys_1_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 52:16]
  wire [15:0] ReApplys_1_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_io_remote_out_ready; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 52:16]
  wire [511:0] ReApplys_1_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 52:16]
  wire [63:0] ReApplys_1_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_io_remote_out_bits_tlast; // @[nf_arm_doce_top_main.scala 52:16]
  wire [3:0] ReApplys_1_io_recv_sync; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_io_recv_sync_phase2; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_io_signal; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_io_signal_ack; // @[nf_arm_doce_top_main.scala 52:16]
  wire [1:0] ReApplys_1_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_1_io_end; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_1_io_packet_size; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_1_io_level; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_1_io_pending_time; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_1_io_pending_parameter; // @[nf_arm_doce_top_main.scala 52:16]
  wire [1:0] ReApplys_1_io_idol_fpga_num; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_clock; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_reset; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 52:16]
  wire [511:0] ReApplys_2_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 52:16]
  wire [15:0] ReApplys_2_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_io_remote_out_ready; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 52:16]
  wire [511:0] ReApplys_2_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 52:16]
  wire [63:0] ReApplys_2_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_io_remote_out_bits_tlast; // @[nf_arm_doce_top_main.scala 52:16]
  wire [3:0] ReApplys_2_io_recv_sync; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_io_recv_sync_phase2; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_io_signal; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_io_signal_ack; // @[nf_arm_doce_top_main.scala 52:16]
  wire [1:0] ReApplys_2_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_2_io_end; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_2_io_packet_size; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_2_io_level; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_2_io_pending_time; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_2_io_pending_parameter; // @[nf_arm_doce_top_main.scala 52:16]
  wire [1:0] ReApplys_2_io_idol_fpga_num; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_clock; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_reset; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 52:16]
  wire [511:0] ReApplys_3_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 52:16]
  wire [15:0] ReApplys_3_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_io_remote_out_ready; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 52:16]
  wire [511:0] ReApplys_3_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 52:16]
  wire [63:0] ReApplys_3_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_io_remote_out_bits_tlast; // @[nf_arm_doce_top_main.scala 52:16]
  wire [3:0] ReApplys_3_io_recv_sync; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_io_recv_sync_phase2; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_io_signal; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_io_signal_ack; // @[nf_arm_doce_top_main.scala 52:16]
  wire [1:0] ReApplys_3_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReApplys_3_io_end; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_3_io_packet_size; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_3_io_level; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_3_io_pending_time; // @[nf_arm_doce_top_main.scala 52:16]
  wire [31:0] ReApplys_3_io_pending_parameter; // @[nf_arm_doce_top_main.scala 52:16]
  wire [1:0] ReApplys_3_io_idol_fpga_num; // @[nf_arm_doce_top_main.scala 52:16]
  wire  ReScatter_clock; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_reset; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_remote_in_w_ready; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_remote_in_w_valid; // @[nf_arm_doce_top_main.scala 54:25]
  wire [511:0] ReScatter_io_remote_in_w_bits_wdata; // @[nf_arm_doce_top_main.scala 54:25]
  wire [63:0] ReScatter_io_remote_in_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 54:25]
  wire [511:0] ReScatter_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 54:25]
  wire [15:0] ReScatter_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_signal; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_start; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_issue_sync; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_issue_sync_phase2_0; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_issue_sync_phase2_1; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_issue_sync_phase2_2; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReScatter_io_issue_sync_phase2_3; // @[nf_arm_doce_top_main.scala 54:25]
  wire [1:0] ReScatter_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 54:25]
  wire [1:0] ReScatter_io_idol_fpga_num; // @[nf_arm_doce_top_main.scala 54:25]
  wire  ReSwitch_clock; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_reset; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_0_ready; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_0_valid; // @[nf_arm_doce_top_main.scala 56:24]
  wire [511:0] ReSwitch_io_xbar_in_0_bits_tdata; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_xbar_in_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_0_bits_tlast; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_1_ready; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_1_valid; // @[nf_arm_doce_top_main.scala 56:24]
  wire [511:0] ReSwitch_io_xbar_in_1_bits_tdata; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_xbar_in_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_1_bits_tlast; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_2_ready; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_2_valid; // @[nf_arm_doce_top_main.scala 56:24]
  wire [511:0] ReSwitch_io_xbar_in_2_bits_tdata; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_xbar_in_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_2_bits_tlast; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_3_ready; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_3_valid; // @[nf_arm_doce_top_main.scala 56:24]
  wire [511:0] ReSwitch_io_xbar_in_3_bits_tdata; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_xbar_in_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_xbar_in_3_bits_tlast; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_remote_out_aw_ready; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_remote_out_aw_valid; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_remote_out_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_remote_out_w_ready; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_remote_out_w_valid; // @[nf_arm_doce_top_main.scala 56:24]
  wire [511:0] ReSwitch_io_remote_out_w_bits_wdata; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_remote_out_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 56:24]
  wire  ReSwitch_io_remote_out_w_bits_wlast; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_level_base_addr_0; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_level_base_addr_1; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_level_base_addr_2; // @[nf_arm_doce_top_main.scala 56:24]
  wire [63:0] ReSwitch_io_level_base_addr_3; // @[nf_arm_doce_top_main.scala 56:24]
  wire [31:0] ReSwitch_io_net_constrain; // @[nf_arm_doce_top_main.scala 56:24]
  reg [31:0] max_size_to_net; // @[nf_arm_doce_top_main.scala 59:32]
  reg [31:0] size_to_net; // @[nf_arm_doce_top_main.scala 61:28]
  wire [31:0] _size_to_net_T_1 = size_to_net + 32'h40; // @[nf_arm_doce_top_main.scala 63:32]
  wire [63:0] _controls_io_traveled_edges_T_1 = Scatters_0_io_traveled_edges + Scatters_1_io_traveled_edges; // @[nf_arm_doce_top_main.scala 119:80]
  wire [63:0] _controls_io_traveled_edges_T_3 = _controls_io_traveled_edges_T_1 + Scatters_2_io_traveled_edges; // @[nf_arm_doce_top_main.scala 119:80]
  wire  _controls_io_signal_ack_T = 32'h0 == controls_io_data_16; // @[nf_arm_doce_top_main.scala 123:41]
  wire  _controls_io_signal_ack_T_1 = ReApplys_0_io_signal_ack | 32'h0 == controls_io_data_16; // @[nf_arm_doce_top_main.scala 123:34]
  wire  _controls_io_signal_ack_T_2 = 32'h1 == controls_io_data_16; // @[nf_arm_doce_top_main.scala 123:41]
  wire  _controls_io_signal_ack_T_3 = ReApplys_1_io_signal_ack | 32'h1 == controls_io_data_16; // @[nf_arm_doce_top_main.scala 123:34]
  wire  _controls_io_signal_ack_T_4 = 32'h2 == controls_io_data_16; // @[nf_arm_doce_top_main.scala 123:41]
  wire  _controls_io_signal_ack_T_5 = ReApplys_2_io_signal_ack | 32'h2 == controls_io_data_16; // @[nf_arm_doce_top_main.scala 123:34]
  wire  _controls_io_signal_ack_T_6 = 32'h3 == controls_io_data_16; // @[nf_arm_doce_top_main.scala 123:41]
  wire  _controls_io_signal_ack_T_7 = ReApplys_3_io_signal_ack | 32'h3 == controls_io_data_16; // @[nf_arm_doce_top_main.scala 123:34]
  wire  _controls_io_signal_ack_T_10 = _controls_io_signal_ack_T_1 & _controls_io_signal_ack_T_3 &
    _controls_io_signal_ack_T_5 & _controls_io_signal_ack_T_7; // @[nf_arm_doce_top_main.scala 124:13]
  wire  _Scatters_0_io_recv_sync_WIRE_1 = Scatters_0_io_issue_sync; // @[nf_arm_doce_top_main.scala 140:32 nf_arm_doce_top_main.scala 140:32]
  wire  _Scatters_0_io_recv_sync_WIRE_0 = ReScatter_io_issue_sync; // @[nf_arm_doce_top_main.scala 140:32 nf_arm_doce_top_main.scala 140:32]
  wire [1:0] Scatters_0_io_recv_sync_lo = {_Scatters_0_io_recv_sync_WIRE_1,_Scatters_0_io_recv_sync_WIRE_0}; // @[nf_arm_doce_top_main.scala 140:103]
  wire  _Scatters_0_io_recv_sync_WIRE_4 = Scatters_3_io_issue_sync; // @[nf_arm_doce_top_main.scala 140:32 nf_arm_doce_top_main.scala 140:32]
  wire  _Scatters_0_io_recv_sync_WIRE_3 = Scatters_2_io_issue_sync; // @[nf_arm_doce_top_main.scala 140:32 nf_arm_doce_top_main.scala 140:32]
  wire [1:0] Scatters_0_io_recv_sync_hi_hi = {_Scatters_0_io_recv_sync_WIRE_4,_Scatters_0_io_recv_sync_WIRE_3}; // @[nf_arm_doce_top_main.scala 140:103]
  wire  _Scatters_0_io_recv_sync_WIRE_2 = Scatters_1_io_issue_sync; // @[nf_arm_doce_top_main.scala 140:32 nf_arm_doce_top_main.scala 140:32]
  wire [2:0] Scatters_0_io_recv_sync_hi = {_Scatters_0_io_recv_sync_WIRE_4,_Scatters_0_io_recv_sync_WIRE_3,
    _Scatters_0_io_recv_sync_WIRE_2}; // @[nf_arm_doce_top_main.scala 140:103]
  wire [1:0] ReApplys_0_io_recv_sync_lo = {_Scatters_0_io_recv_sync_WIRE_2,_Scatters_0_io_recv_sync_WIRE_1}; // @[nf_arm_doce_top_main.scala 150:75]
  controller controls ( // @[nf_arm_doce_top_main.scala 30:24]
    .clock(controls_clock),
    .reset(controls_reset),
    .io_data_0(controls_io_data_0),
    .io_data_1(controls_io_data_1),
    .io_data_2(controls_io_data_2),
    .io_data_3(controls_io_data_3),
    .io_data_4(controls_io_data_4),
    .io_data_7(controls_io_data_7),
    .io_data_16(controls_io_data_16),
    .io_data_17(controls_io_data_17),
    .io_data_18(controls_io_data_18),
    .io_data_19(controls_io_data_19),
    .io_data_20(controls_io_data_20),
    .io_data_21(controls_io_data_21),
    .io_data_22(controls_io_data_22),
    .io_data_23(controls_io_data_23),
    .io_data_24(controls_io_data_24),
    .io_data_25(controls_io_data_25),
    .io_data_26(controls_io_data_26),
    .io_data_27(controls_io_data_27),
    .io_data_28(controls_io_data_28),
    .io_data_29(controls_io_data_29),
    .io_fin_0(controls_io_fin_0),
    .io_fin_1(controls_io_fin_1),
    .io_fin_2(controls_io_fin_2),
    .io_fin_3(controls_io_fin_3),
    .io_fin_4(controls_io_fin_4),
    .io_fin_5(controls_io_fin_5),
    .io_fin_6(controls_io_fin_6),
    .io_fin_7(controls_io_fin_7),
    .io_fin_8(controls_io_fin_8),
    .io_fin_9(controls_io_fin_9),
    .io_fin_10(controls_io_fin_10),
    .io_fin_11(controls_io_fin_11),
    .io_fin_12(controls_io_fin_12),
    .io_fin_13(controls_io_fin_13),
    .io_fin_14(controls_io_fin_14),
    .io_fin_15(controls_io_fin_15),
    .io_fin_16(controls_io_fin_16),
    .io_fin_17(controls_io_fin_17),
    .io_fin_18(controls_io_fin_18),
    .io_fin_19(controls_io_fin_19),
    .io_signal(controls_io_signal),
    .io_start(controls_io_start),
    .io_level(controls_io_level),
    .io_traveled_edges(controls_io_traveled_edges),
    .io_config_awaddr(controls_io_config_awaddr),
    .io_config_awvalid(controls_io_config_awvalid),
    .io_config_awready(controls_io_config_awready),
    .io_config_araddr(controls_io_config_araddr),
    .io_config_arvalid(controls_io_config_arvalid),
    .io_config_arready(controls_io_config_arready),
    .io_config_wdata(controls_io_config_wdata),
    .io_config_wvalid(controls_io_config_wvalid),
    .io_config_wready(controls_io_config_wready),
    .io_config_rdata(controls_io_config_rdata),
    .io_config_rvalid(controls_io_config_rvalid),
    .io_config_rready(controls_io_config_rready),
    .io_config_bvalid(controls_io_config_bvalid),
    .io_config_bready(controls_io_config_bready),
    .io_flush_cache(controls_io_flush_cache),
    .io_flush_cache_end(controls_io_flush_cache_end),
    .io_signal_ack(controls_io_signal_ack)
  );
  multi_port_mc MemController ( // @[nf_arm_doce_top_main.scala 39:29]
    .clock(MemController_clock),
    .reset(MemController_reset),
    .io_cacheable_out_ready(MemController_io_cacheable_out_ready),
    .io_cacheable_out_valid(MemController_io_cacheable_out_valid),
    .io_cacheable_out_bits_tdata(MemController_io_cacheable_out_bits_tdata),
    .io_cacheable_out_bits_tkeep(MemController_io_cacheable_out_bits_tkeep),
    .io_graph_scale(MemController_io_graph_scale),
    .io_start(MemController_io_start),
    .io_signal(MemController_io_signal),
    .io_end(MemController_io_end),
    .io_signal_ack(MemController_io_signal_ack)
  );
  Scatter Applys_0 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_0_clock),
    .reset(Applys_0_reset),
    .io_xbar_in_ready(Applys_0_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_0_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_0_io_xbar_in_bits_tlast),
    .io_end(Applys_0_io_end),
    .io_local_fpga_id(Applys_0_io_local_fpga_id),
    .io_graph_scale(Applys_0_io_graph_scale)
  );
  Scatter_1 Applys_1 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_1_clock),
    .reset(Applys_1_reset),
    .io_xbar_in_ready(Applys_1_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_1_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_1_io_xbar_in_bits_tlast),
    .io_end(Applys_1_io_end),
    .io_local_fpga_id(Applys_1_io_local_fpga_id),
    .io_graph_scale(Applys_1_io_graph_scale)
  );
  Scatter_2 Applys_2 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_2_clock),
    .reset(Applys_2_reset),
    .io_xbar_in_ready(Applys_2_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_2_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_2_io_xbar_in_bits_tlast),
    .io_end(Applys_2_io_end),
    .io_local_fpga_id(Applys_2_io_local_fpga_id),
    .io_graph_scale(Applys_2_io_graph_scale)
  );
  Scatter_3 Applys_3 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_3_clock),
    .reset(Applys_3_reset),
    .io_xbar_in_ready(Applys_3_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_3_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_3_io_xbar_in_bits_tlast),
    .io_end(Applys_3_io_end),
    .io_local_fpga_id(Applys_3_io_local_fpga_id),
    .io_graph_scale(Applys_3_io_graph_scale)
  );
  Scatter_4 Applys_4 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_4_clock),
    .reset(Applys_4_reset),
    .io_xbar_in_ready(Applys_4_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_4_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_4_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_4_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_4_io_xbar_in_bits_tlast),
    .io_end(Applys_4_io_end),
    .io_local_fpga_id(Applys_4_io_local_fpga_id),
    .io_graph_scale(Applys_4_io_graph_scale)
  );
  Scatter_5 Applys_5 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_5_clock),
    .reset(Applys_5_reset),
    .io_xbar_in_ready(Applys_5_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_5_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_5_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_5_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_5_io_xbar_in_bits_tlast),
    .io_end(Applys_5_io_end),
    .io_local_fpga_id(Applys_5_io_local_fpga_id),
    .io_graph_scale(Applys_5_io_graph_scale)
  );
  Scatter_6 Applys_6 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_6_clock),
    .reset(Applys_6_reset),
    .io_xbar_in_ready(Applys_6_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_6_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_6_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_6_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_6_io_xbar_in_bits_tlast),
    .io_end(Applys_6_io_end),
    .io_local_fpga_id(Applys_6_io_local_fpga_id),
    .io_graph_scale(Applys_6_io_graph_scale)
  );
  Scatter_7 Applys_7 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_7_clock),
    .reset(Applys_7_reset),
    .io_xbar_in_ready(Applys_7_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_7_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_7_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_7_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_7_io_xbar_in_bits_tlast),
    .io_end(Applys_7_io_end),
    .io_local_fpga_id(Applys_7_io_local_fpga_id),
    .io_graph_scale(Applys_7_io_graph_scale)
  );
  Scatter_8 Applys_8 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_8_clock),
    .reset(Applys_8_reset),
    .io_xbar_in_ready(Applys_8_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_8_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_8_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_8_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_8_io_xbar_in_bits_tlast),
    .io_end(Applys_8_io_end),
    .io_local_fpga_id(Applys_8_io_local_fpga_id),
    .io_graph_scale(Applys_8_io_graph_scale)
  );
  Scatter_9 Applys_9 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_9_clock),
    .reset(Applys_9_reset),
    .io_xbar_in_ready(Applys_9_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_9_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_9_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_9_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_9_io_xbar_in_bits_tlast),
    .io_end(Applys_9_io_end),
    .io_local_fpga_id(Applys_9_io_local_fpga_id),
    .io_graph_scale(Applys_9_io_graph_scale)
  );
  Scatter_10 Applys_10 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_10_clock),
    .reset(Applys_10_reset),
    .io_xbar_in_ready(Applys_10_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_10_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_10_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_10_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_10_io_xbar_in_bits_tlast),
    .io_end(Applys_10_io_end),
    .io_local_fpga_id(Applys_10_io_local_fpga_id),
    .io_graph_scale(Applys_10_io_graph_scale)
  );
  Scatter_11 Applys_11 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_11_clock),
    .reset(Applys_11_reset),
    .io_xbar_in_ready(Applys_11_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_11_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_11_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_11_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_11_io_xbar_in_bits_tlast),
    .io_end(Applys_11_io_end),
    .io_local_fpga_id(Applys_11_io_local_fpga_id),
    .io_graph_scale(Applys_11_io_graph_scale)
  );
  Scatter_12 Applys_12 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_12_clock),
    .reset(Applys_12_reset),
    .io_xbar_in_ready(Applys_12_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_12_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_12_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_12_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_12_io_xbar_in_bits_tlast),
    .io_end(Applys_12_io_end),
    .io_local_fpga_id(Applys_12_io_local_fpga_id),
    .io_graph_scale(Applys_12_io_graph_scale)
  );
  Scatter_13 Applys_13 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_13_clock),
    .reset(Applys_13_reset),
    .io_xbar_in_ready(Applys_13_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_13_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_13_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_13_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_13_io_xbar_in_bits_tlast),
    .io_end(Applys_13_io_end),
    .io_local_fpga_id(Applys_13_io_local_fpga_id),
    .io_graph_scale(Applys_13_io_graph_scale)
  );
  Scatter_14 Applys_14 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_14_clock),
    .reset(Applys_14_reset),
    .io_xbar_in_ready(Applys_14_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_14_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_14_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_14_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_14_io_xbar_in_bits_tlast),
    .io_end(Applys_14_io_end),
    .io_local_fpga_id(Applys_14_io_local_fpga_id),
    .io_graph_scale(Applys_14_io_graph_scale)
  );
  Scatter_15 Applys_15 ( // @[nf_arm_doce_top_main.scala 42:16]
    .clock(Applys_15_clock),
    .reset(Applys_15_reset),
    .io_xbar_in_ready(Applys_15_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_15_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_15_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_15_io_xbar_in_bits_tkeep),
    .io_xbar_in_bits_tlast(Applys_15_io_xbar_in_bits_tlast),
    .io_end(Applys_15_io_end),
    .io_local_fpga_id(Applys_15_io_local_fpga_id),
    .io_graph_scale(Applys_15_io_graph_scale)
  );
  Gather Gathers ( // @[nf_arm_doce_top_main.scala 44:23]
    .clock(Gathers_clock),
    .reset(Gathers_reset),
    .io_ddr_in_ready(Gathers_io_ddr_in_ready),
    .io_ddr_in_valid(Gathers_io_ddr_in_valid),
    .io_ddr_in_bits_tdata(Gathers_io_ddr_in_bits_tdata),
    .io_ddr_in_bits_tkeep(Gathers_io_ddr_in_bits_tkeep),
    .io_gather_out_0_ready(Gathers_io_gather_out_0_ready),
    .io_gather_out_0_valid(Gathers_io_gather_out_0_valid),
    .io_gather_out_0_bits_tdata(Gathers_io_gather_out_0_bits_tdata),
    .io_gather_out_1_ready(Gathers_io_gather_out_1_ready),
    .io_gather_out_1_valid(Gathers_io_gather_out_1_valid),
    .io_gather_out_1_bits_tdata(Gathers_io_gather_out_1_bits_tdata),
    .io_gather_out_2_ready(Gathers_io_gather_out_2_ready),
    .io_gather_out_2_valid(Gathers_io_gather_out_2_valid),
    .io_gather_out_2_bits_tdata(Gathers_io_gather_out_2_bits_tdata),
    .io_gather_out_3_ready(Gathers_io_gather_out_3_ready),
    .io_gather_out_3_valid(Gathers_io_gather_out_3_valid),
    .io_gather_out_3_bits_tdata(Gathers_io_gather_out_3_bits_tdata)
  );
  Apply LevelCache ( // @[nf_arm_doce_top_main.scala 45:26]
    .io_end(LevelCache_io_end),
    .io_flush(LevelCache_io_flush)
  );
  Broadcast Scatters_0 ( // @[nf_arm_doce_top_main.scala 47:16]
    .clock(Scatters_0_clock),
    .reset(Scatters_0_reset),
    .io_ddr_ar_ready(Scatters_0_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_0_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_0_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_0_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_0_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_0_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_0_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_0_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_0_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_0_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_0_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_0_io_gather_in_ready),
    .io_gather_in_valid(Scatters_0_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_0_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_0_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_0_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_0_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_0_io_xbar_out_bits_tkeep),
    .io_xbar_out_bits_tlast(Scatters_0_io_xbar_out_bits_tlast),
    .io_embedding_base_addr(Scatters_0_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_0_io_edge_base_addr),
    .io_signal(Scatters_0_io_signal),
    .io_traveled_edges(Scatters_0_io_traveled_edges),
    .io_start(Scatters_0_io_start),
    .io_root(Scatters_0_io_root),
    .io_issue_sync(Scatters_0_io_issue_sync),
    .io_recv_sync(Scatters_0_io_recv_sync)
  );
  Broadcast_1 Scatters_1 ( // @[nf_arm_doce_top_main.scala 47:16]
    .clock(Scatters_1_clock),
    .reset(Scatters_1_reset),
    .io_ddr_ar_ready(Scatters_1_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_1_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_1_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_1_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_1_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_1_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_1_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_1_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_1_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_1_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_1_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_1_io_gather_in_ready),
    .io_gather_in_valid(Scatters_1_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_1_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_1_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_1_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_1_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_1_io_xbar_out_bits_tkeep),
    .io_xbar_out_bits_tlast(Scatters_1_io_xbar_out_bits_tlast),
    .io_embedding_base_addr(Scatters_1_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_1_io_edge_base_addr),
    .io_signal(Scatters_1_io_signal),
    .io_traveled_edges(Scatters_1_io_traveled_edges),
    .io_issue_sync(Scatters_1_io_issue_sync),
    .io_recv_sync(Scatters_1_io_recv_sync)
  );
  Broadcast_2 Scatters_2 ( // @[nf_arm_doce_top_main.scala 47:16]
    .clock(Scatters_2_clock),
    .reset(Scatters_2_reset),
    .io_ddr_ar_ready(Scatters_2_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_2_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_2_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_2_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_2_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_2_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_2_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_2_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_2_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_2_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_2_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_2_io_gather_in_ready),
    .io_gather_in_valid(Scatters_2_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_2_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_2_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_2_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_2_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_2_io_xbar_out_bits_tkeep),
    .io_xbar_out_bits_tlast(Scatters_2_io_xbar_out_bits_tlast),
    .io_embedding_base_addr(Scatters_2_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_2_io_edge_base_addr),
    .io_signal(Scatters_2_io_signal),
    .io_traveled_edges(Scatters_2_io_traveled_edges),
    .io_issue_sync(Scatters_2_io_issue_sync),
    .io_recv_sync(Scatters_2_io_recv_sync)
  );
  Broadcast_3 Scatters_3 ( // @[nf_arm_doce_top_main.scala 47:16]
    .clock(Scatters_3_clock),
    .reset(Scatters_3_reset),
    .io_ddr_ar_ready(Scatters_3_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_3_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_3_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_3_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_3_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_3_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_3_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_3_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_3_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_3_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_3_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_3_io_gather_in_ready),
    .io_gather_in_valid(Scatters_3_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_3_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_3_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_3_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_3_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_3_io_xbar_out_bits_tkeep),
    .io_xbar_out_bits_tlast(Scatters_3_io_xbar_out_bits_tlast),
    .io_embedding_base_addr(Scatters_3_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_3_io_edge_base_addr),
    .io_signal(Scatters_3_io_signal),
    .io_traveled_edges(Scatters_3_io_traveled_edges),
    .io_issue_sync(Scatters_3_io_issue_sync),
    .io_recv_sync(Scatters_3_io_recv_sync)
  );
  Remote_xbar Broadcaster ( // @[nf_arm_doce_top_main.scala 50:27]
    .clock(Broadcaster_clock),
    .reset(Broadcaster_reset),
    .io_ddr_in_0_ready(Broadcaster_io_ddr_in_0_ready),
    .io_ddr_in_0_valid(Broadcaster_io_ddr_in_0_valid),
    .io_ddr_in_0_bits_tdata(Broadcaster_io_ddr_in_0_bits_tdata),
    .io_ddr_in_0_bits_tkeep(Broadcaster_io_ddr_in_0_bits_tkeep),
    .io_ddr_in_0_bits_tlast(Broadcaster_io_ddr_in_0_bits_tlast),
    .io_ddr_in_1_ready(Broadcaster_io_ddr_in_1_ready),
    .io_ddr_in_1_valid(Broadcaster_io_ddr_in_1_valid),
    .io_ddr_in_1_bits_tdata(Broadcaster_io_ddr_in_1_bits_tdata),
    .io_ddr_in_1_bits_tkeep(Broadcaster_io_ddr_in_1_bits_tkeep),
    .io_ddr_in_1_bits_tlast(Broadcaster_io_ddr_in_1_bits_tlast),
    .io_ddr_in_2_ready(Broadcaster_io_ddr_in_2_ready),
    .io_ddr_in_2_valid(Broadcaster_io_ddr_in_2_valid),
    .io_ddr_in_2_bits_tdata(Broadcaster_io_ddr_in_2_bits_tdata),
    .io_ddr_in_2_bits_tkeep(Broadcaster_io_ddr_in_2_bits_tkeep),
    .io_ddr_in_2_bits_tlast(Broadcaster_io_ddr_in_2_bits_tlast),
    .io_ddr_in_3_ready(Broadcaster_io_ddr_in_3_ready),
    .io_ddr_in_3_valid(Broadcaster_io_ddr_in_3_valid),
    .io_ddr_in_3_bits_tdata(Broadcaster_io_ddr_in_3_bits_tdata),
    .io_ddr_in_3_bits_tkeep(Broadcaster_io_ddr_in_3_bits_tkeep),
    .io_ddr_in_3_bits_tlast(Broadcaster_io_ddr_in_3_bits_tlast),
    .io_pe_out_0_ready(Broadcaster_io_pe_out_0_ready),
    .io_pe_out_0_valid(Broadcaster_io_pe_out_0_valid),
    .io_pe_out_0_bits_tdata(Broadcaster_io_pe_out_0_bits_tdata),
    .io_pe_out_0_bits_tkeep(Broadcaster_io_pe_out_0_bits_tkeep),
    .io_pe_out_0_bits_tlast(Broadcaster_io_pe_out_0_bits_tlast),
    .io_pe_out_1_ready(Broadcaster_io_pe_out_1_ready),
    .io_pe_out_1_valid(Broadcaster_io_pe_out_1_valid),
    .io_pe_out_1_bits_tdata(Broadcaster_io_pe_out_1_bits_tdata),
    .io_pe_out_1_bits_tkeep(Broadcaster_io_pe_out_1_bits_tkeep),
    .io_pe_out_1_bits_tlast(Broadcaster_io_pe_out_1_bits_tlast),
    .io_pe_out_2_ready(Broadcaster_io_pe_out_2_ready),
    .io_pe_out_2_valid(Broadcaster_io_pe_out_2_valid),
    .io_pe_out_2_bits_tdata(Broadcaster_io_pe_out_2_bits_tdata),
    .io_pe_out_2_bits_tkeep(Broadcaster_io_pe_out_2_bits_tkeep),
    .io_pe_out_2_bits_tlast(Broadcaster_io_pe_out_2_bits_tlast),
    .io_pe_out_3_ready(Broadcaster_io_pe_out_3_ready),
    .io_pe_out_3_valid(Broadcaster_io_pe_out_3_valid),
    .io_pe_out_3_bits_tdata(Broadcaster_io_pe_out_3_bits_tdata),
    .io_pe_out_3_bits_tkeep(Broadcaster_io_pe_out_3_bits_tkeep),
    .io_pe_out_3_bits_tlast(Broadcaster_io_pe_out_3_bits_tlast),
    .io_pe_out_4_ready(Broadcaster_io_pe_out_4_ready),
    .io_pe_out_4_valid(Broadcaster_io_pe_out_4_valid),
    .io_pe_out_4_bits_tdata(Broadcaster_io_pe_out_4_bits_tdata),
    .io_pe_out_4_bits_tkeep(Broadcaster_io_pe_out_4_bits_tkeep),
    .io_pe_out_4_bits_tlast(Broadcaster_io_pe_out_4_bits_tlast),
    .io_pe_out_5_ready(Broadcaster_io_pe_out_5_ready),
    .io_pe_out_5_valid(Broadcaster_io_pe_out_5_valid),
    .io_pe_out_5_bits_tdata(Broadcaster_io_pe_out_5_bits_tdata),
    .io_pe_out_5_bits_tkeep(Broadcaster_io_pe_out_5_bits_tkeep),
    .io_pe_out_5_bits_tlast(Broadcaster_io_pe_out_5_bits_tlast),
    .io_pe_out_6_ready(Broadcaster_io_pe_out_6_ready),
    .io_pe_out_6_valid(Broadcaster_io_pe_out_6_valid),
    .io_pe_out_6_bits_tdata(Broadcaster_io_pe_out_6_bits_tdata),
    .io_pe_out_6_bits_tkeep(Broadcaster_io_pe_out_6_bits_tkeep),
    .io_pe_out_6_bits_tlast(Broadcaster_io_pe_out_6_bits_tlast),
    .io_pe_out_7_ready(Broadcaster_io_pe_out_7_ready),
    .io_pe_out_7_valid(Broadcaster_io_pe_out_7_valid),
    .io_pe_out_7_bits_tdata(Broadcaster_io_pe_out_7_bits_tdata),
    .io_pe_out_7_bits_tkeep(Broadcaster_io_pe_out_7_bits_tkeep),
    .io_pe_out_7_bits_tlast(Broadcaster_io_pe_out_7_bits_tlast),
    .io_pe_out_8_ready(Broadcaster_io_pe_out_8_ready),
    .io_pe_out_8_valid(Broadcaster_io_pe_out_8_valid),
    .io_pe_out_8_bits_tdata(Broadcaster_io_pe_out_8_bits_tdata),
    .io_pe_out_8_bits_tkeep(Broadcaster_io_pe_out_8_bits_tkeep),
    .io_pe_out_8_bits_tlast(Broadcaster_io_pe_out_8_bits_tlast),
    .io_pe_out_9_ready(Broadcaster_io_pe_out_9_ready),
    .io_pe_out_9_valid(Broadcaster_io_pe_out_9_valid),
    .io_pe_out_9_bits_tdata(Broadcaster_io_pe_out_9_bits_tdata),
    .io_pe_out_9_bits_tkeep(Broadcaster_io_pe_out_9_bits_tkeep),
    .io_pe_out_9_bits_tlast(Broadcaster_io_pe_out_9_bits_tlast),
    .io_pe_out_10_ready(Broadcaster_io_pe_out_10_ready),
    .io_pe_out_10_valid(Broadcaster_io_pe_out_10_valid),
    .io_pe_out_10_bits_tdata(Broadcaster_io_pe_out_10_bits_tdata),
    .io_pe_out_10_bits_tkeep(Broadcaster_io_pe_out_10_bits_tkeep),
    .io_pe_out_10_bits_tlast(Broadcaster_io_pe_out_10_bits_tlast),
    .io_pe_out_11_ready(Broadcaster_io_pe_out_11_ready),
    .io_pe_out_11_valid(Broadcaster_io_pe_out_11_valid),
    .io_pe_out_11_bits_tdata(Broadcaster_io_pe_out_11_bits_tdata),
    .io_pe_out_11_bits_tkeep(Broadcaster_io_pe_out_11_bits_tkeep),
    .io_pe_out_11_bits_tlast(Broadcaster_io_pe_out_11_bits_tlast),
    .io_pe_out_12_ready(Broadcaster_io_pe_out_12_ready),
    .io_pe_out_12_valid(Broadcaster_io_pe_out_12_valid),
    .io_pe_out_12_bits_tdata(Broadcaster_io_pe_out_12_bits_tdata),
    .io_pe_out_12_bits_tkeep(Broadcaster_io_pe_out_12_bits_tkeep),
    .io_pe_out_12_bits_tlast(Broadcaster_io_pe_out_12_bits_tlast),
    .io_pe_out_13_ready(Broadcaster_io_pe_out_13_ready),
    .io_pe_out_13_valid(Broadcaster_io_pe_out_13_valid),
    .io_pe_out_13_bits_tdata(Broadcaster_io_pe_out_13_bits_tdata),
    .io_pe_out_13_bits_tkeep(Broadcaster_io_pe_out_13_bits_tkeep),
    .io_pe_out_13_bits_tlast(Broadcaster_io_pe_out_13_bits_tlast),
    .io_pe_out_14_ready(Broadcaster_io_pe_out_14_ready),
    .io_pe_out_14_valid(Broadcaster_io_pe_out_14_valid),
    .io_pe_out_14_bits_tdata(Broadcaster_io_pe_out_14_bits_tdata),
    .io_pe_out_14_bits_tkeep(Broadcaster_io_pe_out_14_bits_tkeep),
    .io_pe_out_14_bits_tlast(Broadcaster_io_pe_out_14_bits_tlast),
    .io_pe_out_15_ready(Broadcaster_io_pe_out_15_ready),
    .io_pe_out_15_valid(Broadcaster_io_pe_out_15_valid),
    .io_pe_out_15_bits_tdata(Broadcaster_io_pe_out_15_bits_tdata),
    .io_pe_out_15_bits_tkeep(Broadcaster_io_pe_out_15_bits_tkeep),
    .io_pe_out_15_bits_tlast(Broadcaster_io_pe_out_15_bits_tlast),
    .io_remote_out_0_ready(Broadcaster_io_remote_out_0_ready),
    .io_remote_out_0_valid(Broadcaster_io_remote_out_0_valid),
    .io_remote_out_0_bits_tdata(Broadcaster_io_remote_out_0_bits_tdata),
    .io_remote_out_0_bits_tkeep(Broadcaster_io_remote_out_0_bits_tkeep),
    .io_remote_out_1_ready(Broadcaster_io_remote_out_1_ready),
    .io_remote_out_1_valid(Broadcaster_io_remote_out_1_valid),
    .io_remote_out_1_bits_tdata(Broadcaster_io_remote_out_1_bits_tdata),
    .io_remote_out_1_bits_tkeep(Broadcaster_io_remote_out_1_bits_tkeep),
    .io_remote_out_2_ready(Broadcaster_io_remote_out_2_ready),
    .io_remote_out_2_valid(Broadcaster_io_remote_out_2_valid),
    .io_remote_out_2_bits_tdata(Broadcaster_io_remote_out_2_bits_tdata),
    .io_remote_out_2_bits_tkeep(Broadcaster_io_remote_out_2_bits_tkeep),
    .io_remote_out_3_ready(Broadcaster_io_remote_out_3_ready),
    .io_remote_out_3_valid(Broadcaster_io_remote_out_3_valid),
    .io_remote_out_3_bits_tdata(Broadcaster_io_remote_out_3_bits_tdata),
    .io_remote_out_3_bits_tkeep(Broadcaster_io_remote_out_3_bits_tkeep),
    .io_remote_in_ready(Broadcaster_io_remote_in_ready),
    .io_remote_in_valid(Broadcaster_io_remote_in_valid),
    .io_remote_in_bits_tdata(Broadcaster_io_remote_in_bits_tdata),
    .io_remote_in_bits_tkeep(Broadcaster_io_remote_in_bits_tkeep),
    .io_local_fpga_id(Broadcaster_io_local_fpga_id),
    .io_flush(Broadcaster_io_flush),
    .io_signal(Broadcaster_io_signal)
  );
  Remote_Apply ReApplys_0 ( // @[nf_arm_doce_top_main.scala 52:16]
    .clock(ReApplys_0_clock),
    .reset(ReApplys_0_reset),
    .io_xbar_in_ready(ReApplys_0_io_xbar_in_ready),
    .io_xbar_in_valid(ReApplys_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(ReApplys_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(ReApplys_0_io_xbar_in_bits_tkeep),
    .io_remote_out_ready(ReApplys_0_io_remote_out_ready),
    .io_remote_out_valid(ReApplys_0_io_remote_out_valid),
    .io_remote_out_bits_tdata(ReApplys_0_io_remote_out_bits_tdata),
    .io_remote_out_bits_tkeep(ReApplys_0_io_remote_out_bits_tkeep),
    .io_remote_out_bits_tlast(ReApplys_0_io_remote_out_bits_tlast),
    .io_recv_sync(ReApplys_0_io_recv_sync),
    .io_recv_sync_phase2(ReApplys_0_io_recv_sync_phase2),
    .io_signal(ReApplys_0_io_signal),
    .io_signal_ack(ReApplys_0_io_signal_ack),
    .io_local_fpga_id(ReApplys_0_io_local_fpga_id),
    .io_end(ReApplys_0_io_end),
    .io_packet_size(ReApplys_0_io_packet_size),
    .io_level(ReApplys_0_io_level),
    .io_pending_time(ReApplys_0_io_pending_time),
    .io_pending_parameter(ReApplys_0_io_pending_parameter),
    .io_idol_fpga_num(ReApplys_0_io_idol_fpga_num)
  );
  Remote_Apply_1 ReApplys_1 ( // @[nf_arm_doce_top_main.scala 52:16]
    .clock(ReApplys_1_clock),
    .reset(ReApplys_1_reset),
    .io_xbar_in_ready(ReApplys_1_io_xbar_in_ready),
    .io_xbar_in_valid(ReApplys_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(ReApplys_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(ReApplys_1_io_xbar_in_bits_tkeep),
    .io_remote_out_ready(ReApplys_1_io_remote_out_ready),
    .io_remote_out_valid(ReApplys_1_io_remote_out_valid),
    .io_remote_out_bits_tdata(ReApplys_1_io_remote_out_bits_tdata),
    .io_remote_out_bits_tkeep(ReApplys_1_io_remote_out_bits_tkeep),
    .io_remote_out_bits_tlast(ReApplys_1_io_remote_out_bits_tlast),
    .io_recv_sync(ReApplys_1_io_recv_sync),
    .io_recv_sync_phase2(ReApplys_1_io_recv_sync_phase2),
    .io_signal(ReApplys_1_io_signal),
    .io_signal_ack(ReApplys_1_io_signal_ack),
    .io_local_fpga_id(ReApplys_1_io_local_fpga_id),
    .io_end(ReApplys_1_io_end),
    .io_packet_size(ReApplys_1_io_packet_size),
    .io_level(ReApplys_1_io_level),
    .io_pending_time(ReApplys_1_io_pending_time),
    .io_pending_parameter(ReApplys_1_io_pending_parameter),
    .io_idol_fpga_num(ReApplys_1_io_idol_fpga_num)
  );
  Remote_Apply_2 ReApplys_2 ( // @[nf_arm_doce_top_main.scala 52:16]
    .clock(ReApplys_2_clock),
    .reset(ReApplys_2_reset),
    .io_xbar_in_ready(ReApplys_2_io_xbar_in_ready),
    .io_xbar_in_valid(ReApplys_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(ReApplys_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(ReApplys_2_io_xbar_in_bits_tkeep),
    .io_remote_out_ready(ReApplys_2_io_remote_out_ready),
    .io_remote_out_valid(ReApplys_2_io_remote_out_valid),
    .io_remote_out_bits_tdata(ReApplys_2_io_remote_out_bits_tdata),
    .io_remote_out_bits_tkeep(ReApplys_2_io_remote_out_bits_tkeep),
    .io_remote_out_bits_tlast(ReApplys_2_io_remote_out_bits_tlast),
    .io_recv_sync(ReApplys_2_io_recv_sync),
    .io_recv_sync_phase2(ReApplys_2_io_recv_sync_phase2),
    .io_signal(ReApplys_2_io_signal),
    .io_signal_ack(ReApplys_2_io_signal_ack),
    .io_local_fpga_id(ReApplys_2_io_local_fpga_id),
    .io_end(ReApplys_2_io_end),
    .io_packet_size(ReApplys_2_io_packet_size),
    .io_level(ReApplys_2_io_level),
    .io_pending_time(ReApplys_2_io_pending_time),
    .io_pending_parameter(ReApplys_2_io_pending_parameter),
    .io_idol_fpga_num(ReApplys_2_io_idol_fpga_num)
  );
  Remote_Apply_3 ReApplys_3 ( // @[nf_arm_doce_top_main.scala 52:16]
    .clock(ReApplys_3_clock),
    .reset(ReApplys_3_reset),
    .io_xbar_in_ready(ReApplys_3_io_xbar_in_ready),
    .io_xbar_in_valid(ReApplys_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(ReApplys_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(ReApplys_3_io_xbar_in_bits_tkeep),
    .io_remote_out_ready(ReApplys_3_io_remote_out_ready),
    .io_remote_out_valid(ReApplys_3_io_remote_out_valid),
    .io_remote_out_bits_tdata(ReApplys_3_io_remote_out_bits_tdata),
    .io_remote_out_bits_tkeep(ReApplys_3_io_remote_out_bits_tkeep),
    .io_remote_out_bits_tlast(ReApplys_3_io_remote_out_bits_tlast),
    .io_recv_sync(ReApplys_3_io_recv_sync),
    .io_recv_sync_phase2(ReApplys_3_io_recv_sync_phase2),
    .io_signal(ReApplys_3_io_signal),
    .io_signal_ack(ReApplys_3_io_signal_ack),
    .io_local_fpga_id(ReApplys_3_io_local_fpga_id),
    .io_end(ReApplys_3_io_end),
    .io_packet_size(ReApplys_3_io_packet_size),
    .io_level(ReApplys_3_io_level),
    .io_pending_time(ReApplys_3_io_pending_time),
    .io_pending_parameter(ReApplys_3_io_pending_parameter),
    .io_idol_fpga_num(ReApplys_3_io_idol_fpga_num)
  );
  Remote_Scatter ReScatter ( // @[nf_arm_doce_top_main.scala 54:25]
    .clock(ReScatter_clock),
    .reset(ReScatter_reset),
    .io_remote_in_w_ready(ReScatter_io_remote_in_w_ready),
    .io_remote_in_w_valid(ReScatter_io_remote_in_w_valid),
    .io_remote_in_w_bits_wdata(ReScatter_io_remote_in_w_bits_wdata),
    .io_remote_in_w_bits_wstrb(ReScatter_io_remote_in_w_bits_wstrb),
    .io_xbar_out_ready(ReScatter_io_xbar_out_ready),
    .io_xbar_out_valid(ReScatter_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(ReScatter_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(ReScatter_io_xbar_out_bits_tkeep),
    .io_signal(ReScatter_io_signal),
    .io_start(ReScatter_io_start),
    .io_issue_sync(ReScatter_io_issue_sync),
    .io_issue_sync_phase2_0(ReScatter_io_issue_sync_phase2_0),
    .io_issue_sync_phase2_1(ReScatter_io_issue_sync_phase2_1),
    .io_issue_sync_phase2_2(ReScatter_io_issue_sync_phase2_2),
    .io_issue_sync_phase2_3(ReScatter_io_issue_sync_phase2_3),
    .io_local_fpga_id(ReScatter_io_local_fpga_id),
    .io_idol_fpga_num(ReScatter_io_idol_fpga_num)
  );
  axis_to_axi ReSwitch ( // @[nf_arm_doce_top_main.scala 56:24]
    .clock(ReSwitch_clock),
    .reset(ReSwitch_reset),
    .io_xbar_in_0_ready(ReSwitch_io_xbar_in_0_ready),
    .io_xbar_in_0_valid(ReSwitch_io_xbar_in_0_valid),
    .io_xbar_in_0_bits_tdata(ReSwitch_io_xbar_in_0_bits_tdata),
    .io_xbar_in_0_bits_tkeep(ReSwitch_io_xbar_in_0_bits_tkeep),
    .io_xbar_in_0_bits_tlast(ReSwitch_io_xbar_in_0_bits_tlast),
    .io_xbar_in_1_ready(ReSwitch_io_xbar_in_1_ready),
    .io_xbar_in_1_valid(ReSwitch_io_xbar_in_1_valid),
    .io_xbar_in_1_bits_tdata(ReSwitch_io_xbar_in_1_bits_tdata),
    .io_xbar_in_1_bits_tkeep(ReSwitch_io_xbar_in_1_bits_tkeep),
    .io_xbar_in_1_bits_tlast(ReSwitch_io_xbar_in_1_bits_tlast),
    .io_xbar_in_2_ready(ReSwitch_io_xbar_in_2_ready),
    .io_xbar_in_2_valid(ReSwitch_io_xbar_in_2_valid),
    .io_xbar_in_2_bits_tdata(ReSwitch_io_xbar_in_2_bits_tdata),
    .io_xbar_in_2_bits_tkeep(ReSwitch_io_xbar_in_2_bits_tkeep),
    .io_xbar_in_2_bits_tlast(ReSwitch_io_xbar_in_2_bits_tlast),
    .io_xbar_in_3_ready(ReSwitch_io_xbar_in_3_ready),
    .io_xbar_in_3_valid(ReSwitch_io_xbar_in_3_valid),
    .io_xbar_in_3_bits_tdata(ReSwitch_io_xbar_in_3_bits_tdata),
    .io_xbar_in_3_bits_tkeep(ReSwitch_io_xbar_in_3_bits_tkeep),
    .io_xbar_in_3_bits_tlast(ReSwitch_io_xbar_in_3_bits_tlast),
    .io_remote_out_aw_ready(ReSwitch_io_remote_out_aw_ready),
    .io_remote_out_aw_valid(ReSwitch_io_remote_out_aw_valid),
    .io_remote_out_aw_bits_awaddr(ReSwitch_io_remote_out_aw_bits_awaddr),
    .io_remote_out_w_ready(ReSwitch_io_remote_out_w_ready),
    .io_remote_out_w_valid(ReSwitch_io_remote_out_w_valid),
    .io_remote_out_w_bits_wdata(ReSwitch_io_remote_out_w_bits_wdata),
    .io_remote_out_w_bits_wstrb(ReSwitch_io_remote_out_w_bits_wstrb),
    .io_remote_out_w_bits_wlast(ReSwitch_io_remote_out_w_bits_wlast),
    .io_level_base_addr_0(ReSwitch_io_level_base_addr_0),
    .io_level_base_addr_1(ReSwitch_io_level_base_addr_1),
    .io_level_base_addr_2(ReSwitch_io_level_base_addr_2),
    .io_level_base_addr_3(ReSwitch_io_level_base_addr_3),
    .io_net_constrain(ReSwitch_io_net_constrain)
  );
  assign io_config_awready = controls_io_config_awready; // @[nf_arm_doce_top_main.scala 118:22]
  assign io_config_arready = controls_io_config_arready; // @[nf_arm_doce_top_main.scala 118:22]
  assign io_config_wready = controls_io_config_wready; // @[nf_arm_doce_top_main.scala 118:22]
  assign io_config_rdata = controls_io_config_rdata; // @[nf_arm_doce_top_main.scala 118:22]
  assign io_config_rresp = 2'h0; // @[nf_arm_doce_top_main.scala 118:22]
  assign io_config_rvalid = controls_io_config_rvalid; // @[nf_arm_doce_top_main.scala 118:22]
  assign io_config_bresp = 2'h0; // @[nf_arm_doce_top_main.scala 118:22]
  assign io_config_bvalid = controls_io_config_bvalid; // @[nf_arm_doce_top_main.scala 118:22]
  assign io_PLmemory_0_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_aw_bits_awid = 7'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_ar_valid = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_ar_bits_araddr = 64'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_ar_bits_arid = 7'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_ar_bits_arlen = 8'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_ar_bits_arsize = 3'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_ar_bits_arburst = 2'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_w_bits_wdata = 512'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_w_bits_wstrb = 64'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_w_bits_wlast = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_r_ready = 1'h1; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_0_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_aw_bits_awid = 7'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_ar_valid = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_ar_bits_araddr = 64'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_ar_bits_arid = 7'h40; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_ar_bits_arlen = 8'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_ar_bits_arsize = 3'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_ar_bits_arburst = 2'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_w_bits_wdata = 512'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_w_bits_wstrb = 64'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_w_bits_wlast = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_r_ready = 1'h0; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PLmemory_1_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 71:15]
  assign io_PSmemory_0_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 108:18]
  assign io_PSmemory_0_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_0_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 52:10]
  assign io_PSmemory_0_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 53:11]
  assign io_PSmemory_0_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 54:12]
  assign io_PSmemory_0_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 55:13]
  assign io_PSmemory_0_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 56:12]
  assign io_PSmemory_0_ar_valid = Scatters_0_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_0_ar_bits_araddr = Scatters_0_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_0_ar_bits_arid = Scatters_0_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_0_ar_bits_arlen = Scatters_0_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_0_ar_bits_arsize = Scatters_0_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_0_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_0_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_0_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 110:17]
  assign io_PSmemory_0_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 66:11]
  assign io_PSmemory_0_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 67:11]
  assign io_PSmemory_0_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 68:11]
  assign io_PSmemory_0_r_ready = Scatters_0_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 80:18]
  assign io_PSmemory_0_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 106:17]
  assign io_PSmemory_1_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 108:18]
  assign io_PSmemory_1_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_1_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 52:10]
  assign io_PSmemory_1_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 53:11]
  assign io_PSmemory_1_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 54:12]
  assign io_PSmemory_1_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 55:13]
  assign io_PSmemory_1_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 56:12]
  assign io_PSmemory_1_ar_valid = Scatters_1_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_1_ar_bits_araddr = Scatters_1_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_1_ar_bits_arid = Scatters_1_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_1_ar_bits_arlen = Scatters_1_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_1_ar_bits_arsize = Scatters_1_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_1_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_1_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_1_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 110:17]
  assign io_PSmemory_1_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 66:11]
  assign io_PSmemory_1_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 67:11]
  assign io_PSmemory_1_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 68:11]
  assign io_PSmemory_1_r_ready = Scatters_1_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 80:18]
  assign io_PSmemory_1_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 106:17]
  assign io_PSmemory_2_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 108:18]
  assign io_PSmemory_2_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_2_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 52:10]
  assign io_PSmemory_2_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 53:11]
  assign io_PSmemory_2_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 54:12]
  assign io_PSmemory_2_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 55:13]
  assign io_PSmemory_2_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 56:12]
  assign io_PSmemory_2_ar_valid = Scatters_2_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_2_ar_bits_araddr = Scatters_2_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_2_ar_bits_arid = Scatters_2_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_2_ar_bits_arlen = Scatters_2_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_2_ar_bits_arsize = Scatters_2_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_2_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_2_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_2_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 110:17]
  assign io_PSmemory_2_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 66:11]
  assign io_PSmemory_2_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 67:11]
  assign io_PSmemory_2_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 68:11]
  assign io_PSmemory_2_r_ready = Scatters_2_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 80:18]
  assign io_PSmemory_2_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 106:17]
  assign io_PSmemory_3_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 108:18]
  assign io_PSmemory_3_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_3_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 52:10]
  assign io_PSmemory_3_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 53:11]
  assign io_PSmemory_3_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 54:12]
  assign io_PSmemory_3_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 55:13]
  assign io_PSmemory_3_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 56:12]
  assign io_PSmemory_3_ar_valid = Scatters_3_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_3_ar_bits_araddr = Scatters_3_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_3_ar_bits_arid = Scatters_3_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_3_ar_bits_arlen = Scatters_3_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_3_ar_bits_arsize = Scatters_3_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_3_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_3_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 81:19]
  assign io_PSmemory_3_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 110:17]
  assign io_PSmemory_3_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 66:11]
  assign io_PSmemory_3_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 67:11]
  assign io_PSmemory_3_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 68:11]
  assign io_PSmemory_3_r_ready = Scatters_3_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 80:18]
  assign io_PSmemory_3_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 106:17]
  assign io_Re_memory_out_aw_valid = ReSwitch_io_remote_out_aw_valid; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_aw_bits_awaddr = ReSwitch_io_remote_out_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_aw_bits_awid = 6'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_aw_bits_awsize = 3'h6; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_ar_valid = 1'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_ar_bits_araddr = 64'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_ar_bits_arid = 6'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_ar_bits_arlen = 8'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_ar_bits_arsize = 3'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_ar_bits_arburst = 2'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_w_valid = ReSwitch_io_remote_out_w_valid; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_w_bits_wdata = ReSwitch_io_remote_out_w_bits_wdata; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_w_bits_wstrb = ReSwitch_io_remote_out_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_w_bits_wlast = ReSwitch_io_remote_out_w_bits_wlast; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_r_ready = 1'h1; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_out_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 101:20]
  assign io_Re_memory_in_aw_ready = 1'h1; // @[nf_arm_doce_top_main.scala 94:26]
  assign io_Re_memory_in_ar_ready = 1'h0; // @[nf_arm_doce_top_main.scala 94:26]
  assign io_Re_memory_in_w_ready = ReScatter_io_remote_in_w_ready; // @[nf_arm_doce_top_main.scala 94:26]
  assign io_Re_memory_in_r_valid = 1'h0; // @[nf_arm_doce_top_main.scala 94:26]
  assign io_Re_memory_in_r_bits_rdata = 512'h0; // @[nf_arm_doce_top_main.scala 94:26]
  assign io_Re_memory_in_r_bits_rid = 10'h0; // @[nf_arm_doce_top_main.scala 94:26]
  assign io_Re_memory_in_r_bits_rlast = 1'h0; // @[nf_arm_doce_top_main.scala 94:26]
  assign io_Re_memory_in_b_valid = 1'h0; // @[nf_arm_doce_top_main.scala 94:26]
  assign io_Re_memory_in_b_bits_bresp = 2'h0; // @[nf_arm_doce_top_main.scala 94:26]
  assign io_Re_memory_in_b_bits_bid = 10'h0; // @[nf_arm_doce_top_main.scala 94:26]
  assign controls_clock = clock;
  assign controls_reset = reset;
  assign controls_io_fin_0 = Applys_0_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_1 = Applys_1_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_2 = Applys_2_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_3 = Applys_3_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_4 = Applys_4_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_5 = Applys_5_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_6 = Applys_6_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_7 = Applys_7_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_8 = Applys_8_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_9 = Applys_9_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_10 = Applys_10_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_11 = Applys_11_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_12 = Applys_12_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_13 = Applys_13_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_14 = Applys_14_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_15 = Applys_15_io_end; // @[nf_arm_doce_top_main.scala 89:26]
  assign controls_io_fin_16 = ReApplys_0_io_end | _controls_io_signal_ack_T; // @[nf_arm_doce_top_main.scala 149:41]
  assign controls_io_fin_17 = ReApplys_1_io_end | _controls_io_signal_ack_T_2; // @[nf_arm_doce_top_main.scala 149:41]
  assign controls_io_fin_18 = ReApplys_2_io_end | _controls_io_signal_ack_T_4; // @[nf_arm_doce_top_main.scala 149:41]
  assign controls_io_fin_19 = ReApplys_3_io_end | _controls_io_signal_ack_T_6; // @[nf_arm_doce_top_main.scala 149:41]
  assign controls_io_traveled_edges = _controls_io_traveled_edges_T_3 + Scatters_3_io_traveled_edges; // @[nf_arm_doce_top_main.scala 119:80]
  assign controls_io_config_awaddr = io_config_awaddr; // @[nf_arm_doce_top_main.scala 118:22]
  assign controls_io_config_awvalid = io_config_awvalid; // @[nf_arm_doce_top_main.scala 118:22]
  assign controls_io_config_araddr = io_config_araddr; // @[nf_arm_doce_top_main.scala 118:22]
  assign controls_io_config_arvalid = io_config_arvalid; // @[nf_arm_doce_top_main.scala 118:22]
  assign controls_io_config_wdata = io_config_wdata; // @[nf_arm_doce_top_main.scala 118:22]
  assign controls_io_config_wvalid = io_config_wvalid; // @[nf_arm_doce_top_main.scala 118:22]
  assign controls_io_config_rready = io_config_rready; // @[nf_arm_doce_top_main.scala 118:22]
  assign controls_io_config_bready = io_config_bready; // @[nf_arm_doce_top_main.scala 118:22]
  assign controls_io_flush_cache_end = LevelCache_io_end; // @[nf_arm_doce_top_main.scala 121:31]
  assign controls_io_signal_ack = MemController_io_signal_ack & _controls_io_signal_ack_T_10; // @[nf_arm_doce_top_main.scala 122:57]
  assign MemController_clock = clock;
  assign MemController_reset = reset;
  assign MemController_io_cacheable_out_ready = Gathers_io_ddr_in_ready; // @[nf_arm_doce_top_main.scala 72:21]
  assign MemController_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 143:32]
  assign MemController_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 145:26]
  assign MemController_io_signal = controls_io_signal & controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 144:49]
  assign MemController_io_end = controls_io_data_0[1]; // @[nf_arm_doce_top_main.scala 146:46]
  assign Applys_0_clock = clock;
  assign Applys_0_reset = reset;
  assign Applys_0_io_xbar_in_valid = Broadcaster_io_pe_out_0_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_0_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_0_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_0_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_0_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_0_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_0_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_1_clock = clock;
  assign Applys_1_reset = reset;
  assign Applys_1_io_xbar_in_valid = Broadcaster_io_pe_out_1_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_1_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_1_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_1_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_1_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_1_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_1_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_2_clock = clock;
  assign Applys_2_reset = reset;
  assign Applys_2_io_xbar_in_valid = Broadcaster_io_pe_out_2_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_2_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_2_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_2_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_2_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_2_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_2_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_3_clock = clock;
  assign Applys_3_reset = reset;
  assign Applys_3_io_xbar_in_valid = Broadcaster_io_pe_out_3_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_3_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_3_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_3_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_3_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_3_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_3_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_4_clock = clock;
  assign Applys_4_reset = reset;
  assign Applys_4_io_xbar_in_valid = Broadcaster_io_pe_out_4_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_4_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_4_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_4_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_4_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_4_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_4_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_4_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_5_clock = clock;
  assign Applys_5_reset = reset;
  assign Applys_5_io_xbar_in_valid = Broadcaster_io_pe_out_5_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_5_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_5_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_5_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_5_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_5_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_5_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_5_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_5_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_6_clock = clock;
  assign Applys_6_reset = reset;
  assign Applys_6_io_xbar_in_valid = Broadcaster_io_pe_out_6_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_6_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_6_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_6_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_6_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_6_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_6_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_6_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_6_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_7_clock = clock;
  assign Applys_7_reset = reset;
  assign Applys_7_io_xbar_in_valid = Broadcaster_io_pe_out_7_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_7_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_7_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_7_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_7_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_7_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_7_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_7_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_7_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_8_clock = clock;
  assign Applys_8_reset = reset;
  assign Applys_8_io_xbar_in_valid = Broadcaster_io_pe_out_8_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_8_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_8_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_8_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_8_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_8_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_8_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_8_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_8_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_9_clock = clock;
  assign Applys_9_reset = reset;
  assign Applys_9_io_xbar_in_valid = Broadcaster_io_pe_out_9_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_9_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_9_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_9_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_9_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_9_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_9_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_9_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_9_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_10_clock = clock;
  assign Applys_10_reset = reset;
  assign Applys_10_io_xbar_in_valid = Broadcaster_io_pe_out_10_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_10_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_10_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_10_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_10_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_10_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_10_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_10_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_10_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_11_clock = clock;
  assign Applys_11_reset = reset;
  assign Applys_11_io_xbar_in_valid = Broadcaster_io_pe_out_11_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_11_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_11_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_11_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_11_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_11_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_11_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_11_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_11_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_12_clock = clock;
  assign Applys_12_reset = reset;
  assign Applys_12_io_xbar_in_valid = Broadcaster_io_pe_out_12_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_12_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_12_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_12_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_12_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_12_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_12_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_12_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_12_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_13_clock = clock;
  assign Applys_13_reset = reset;
  assign Applys_13_io_xbar_in_valid = Broadcaster_io_pe_out_13_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_13_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_13_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_13_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_13_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_13_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_13_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_13_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_13_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_14_clock = clock;
  assign Applys_14_reset = reset;
  assign Applys_14_io_xbar_in_valid = Broadcaster_io_pe_out_14_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_14_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_14_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_14_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_14_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_14_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_14_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_14_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_14_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Applys_15_clock = clock;
  assign Applys_15_reset = reset;
  assign Applys_15_io_xbar_in_valid = Broadcaster_io_pe_out_15_valid; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_15_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_15_bits_tdata; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_15_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_15_bits_tkeep; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_15_io_xbar_in_bits_tlast = Broadcaster_io_pe_out_15_bits_tlast; // @[nf_arm_doce_top_main.scala 87:21]
  assign Applys_15_io_local_fpga_id = controls_io_data_16[2:0]; // @[nf_arm_doce_top_main.scala 162:38]
  assign Applys_15_io_graph_scale = controls_io_data_29; // @[nf_arm_doce_top_main.scala 90:25]
  assign Gathers_clock = clock;
  assign Gathers_reset = reset;
  assign Gathers_io_ddr_in_valid = MemController_io_cacheable_out_valid; // @[nf_arm_doce_top_main.scala 72:21]
  assign Gathers_io_ddr_in_bits_tdata = MemController_io_cacheable_out_bits_tdata; // @[nf_arm_doce_top_main.scala 72:21]
  assign Gathers_io_ddr_in_bits_tkeep = MemController_io_cacheable_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 72:21]
  assign Gathers_io_gather_out_0_ready = Scatters_0_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 79:22]
  assign Gathers_io_gather_out_1_ready = Scatters_1_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 79:22]
  assign Gathers_io_gather_out_2_ready = Scatters_2_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 79:22]
  assign Gathers_io_gather_out_3_ready = Scatters_3_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 79:22]
  assign LevelCache_io_flush = controls_io_flush_cache; // @[nf_arm_doce_top_main.scala 126:23]
  assign Scatters_0_clock = clock;
  assign Scatters_0_reset = reset;
  assign Scatters_0_io_ddr_ar_ready = io_PSmemory_0_ar_ready; // @[nf_arm_doce_top_main.scala 81:19]
  assign Scatters_0_io_ddr_r_valid = io_PSmemory_0_r_valid; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_0_io_ddr_r_bits_rdata = io_PSmemory_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_0_io_ddr_r_bits_rid = io_PSmemory_0_r_bits_rid; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_0_io_ddr_r_bits_rlast = io_PSmemory_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_0_io_gather_in_valid = Gathers_io_gather_out_0_valid; // @[nf_arm_doce_top_main.scala 79:22]
  assign Scatters_0_io_gather_in_bits_tdata = Gathers_io_gather_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 79:22]
  assign Scatters_0_io_xbar_out_ready = Broadcaster_io_ddr_in_0_ready; // @[nf_arm_doce_top_main.scala 82:32]
  assign Scatters_0_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_0_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_0_io_signal = controls_io_signal & controls_io_signal_ack | controls_io_start; // @[nf_arm_doce_top_main.scala 132:69]
  assign Scatters_0_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 136:20]
  assign Scatters_0_io_root = controls_io_data_7; // @[nf_arm_doce_top_main.scala 131:17]
  assign Scatters_0_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 140:103]
  assign Scatters_1_clock = clock;
  assign Scatters_1_reset = reset;
  assign Scatters_1_io_ddr_ar_ready = io_PSmemory_1_ar_ready; // @[nf_arm_doce_top_main.scala 81:19]
  assign Scatters_1_io_ddr_r_valid = io_PSmemory_1_r_valid; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_1_io_ddr_r_bits_rdata = io_PSmemory_1_r_bits_rdata; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_1_io_ddr_r_bits_rid = io_PSmemory_1_r_bits_rid; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_1_io_ddr_r_bits_rlast = io_PSmemory_1_r_bits_rlast; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_1_io_gather_in_valid = Gathers_io_gather_out_1_valid; // @[nf_arm_doce_top_main.scala 79:22]
  assign Scatters_1_io_gather_in_bits_tdata = Gathers_io_gather_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 79:22]
  assign Scatters_1_io_xbar_out_ready = Broadcaster_io_ddr_in_1_ready; // @[nf_arm_doce_top_main.scala 82:32]
  assign Scatters_1_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_1_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_1_io_signal = controls_io_signal & controls_io_signal_ack | controls_io_start; // @[nf_arm_doce_top_main.scala 132:69]
  assign Scatters_1_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 140:103]
  assign Scatters_2_clock = clock;
  assign Scatters_2_reset = reset;
  assign Scatters_2_io_ddr_ar_ready = io_PSmemory_2_ar_ready; // @[nf_arm_doce_top_main.scala 81:19]
  assign Scatters_2_io_ddr_r_valid = io_PSmemory_2_r_valid; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_2_io_ddr_r_bits_rdata = io_PSmemory_2_r_bits_rdata; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_2_io_ddr_r_bits_rid = io_PSmemory_2_r_bits_rid; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_2_io_ddr_r_bits_rlast = io_PSmemory_2_r_bits_rlast; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_2_io_gather_in_valid = Gathers_io_gather_out_2_valid; // @[nf_arm_doce_top_main.scala 79:22]
  assign Scatters_2_io_gather_in_bits_tdata = Gathers_io_gather_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 79:22]
  assign Scatters_2_io_xbar_out_ready = Broadcaster_io_ddr_in_2_ready; // @[nf_arm_doce_top_main.scala 82:32]
  assign Scatters_2_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_2_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_2_io_signal = controls_io_signal & controls_io_signal_ack | controls_io_start; // @[nf_arm_doce_top_main.scala 132:69]
  assign Scatters_2_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 140:103]
  assign Scatters_3_clock = clock;
  assign Scatters_3_reset = reset;
  assign Scatters_3_io_ddr_ar_ready = io_PSmemory_3_ar_ready; // @[nf_arm_doce_top_main.scala 81:19]
  assign Scatters_3_io_ddr_r_valid = io_PSmemory_3_r_valid; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_3_io_ddr_r_bits_rdata = io_PSmemory_3_r_bits_rdata; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_3_io_ddr_r_bits_rid = io_PSmemory_3_r_bits_rid; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_3_io_ddr_r_bits_rlast = io_PSmemory_3_r_bits_rlast; // @[nf_arm_doce_top_main.scala 80:18]
  assign Scatters_3_io_gather_in_valid = Gathers_io_gather_out_3_valid; // @[nf_arm_doce_top_main.scala 79:22]
  assign Scatters_3_io_gather_in_bits_tdata = Gathers_io_gather_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 79:22]
  assign Scatters_3_io_xbar_out_ready = Broadcaster_io_ddr_in_3_ready; // @[nf_arm_doce_top_main.scala 82:32]
  assign Scatters_3_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_3_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_3_io_signal = controls_io_signal & controls_io_signal_ack | controls_io_start; // @[nf_arm_doce_top_main.scala 132:69]
  assign Scatters_3_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 140:103]
  assign Broadcaster_clock = clock;
  assign Broadcaster_reset = reset;
  assign Broadcaster_io_ddr_in_0_valid = Scatters_0_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_0_bits_tdata = Scatters_0_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_0_bits_tkeep = Scatters_0_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_0_bits_tlast = Scatters_0_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_1_valid = Scatters_1_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_1_bits_tdata = Scatters_1_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_1_bits_tkeep = Scatters_1_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_1_bits_tlast = Scatters_1_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_2_valid = Scatters_2_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_2_bits_tdata = Scatters_2_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_2_bits_tkeep = Scatters_2_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_2_bits_tlast = Scatters_2_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_3_valid = Scatters_3_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_3_bits_tdata = Scatters_3_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_3_bits_tkeep = Scatters_3_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_ddr_in_3_bits_tlast = Scatters_3_io_xbar_out_bits_tlast; // @[nf_arm_doce_top_main.scala 82:32]
  assign Broadcaster_io_pe_out_0_ready = Applys_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_1_ready = Applys_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_2_ready = Applys_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_3_ready = Applys_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_4_ready = Applys_4_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_5_ready = Applys_5_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_6_ready = Applys_6_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_7_ready = Applys_7_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_8_ready = Applys_8_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_9_ready = Applys_9_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_10_ready = Applys_10_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_11_ready = Applys_11_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_12_ready = Applys_12_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_13_ready = Applys_13_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_14_ready = Applys_14_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_pe_out_15_ready = Applys_15_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 87:21]
  assign Broadcaster_io_remote_out_0_ready = ReApplys_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 97:20]
  assign Broadcaster_io_remote_out_1_ready = ReApplys_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 97:20]
  assign Broadcaster_io_remote_out_2_ready = ReApplys_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 97:20]
  assign Broadcaster_io_remote_out_3_ready = ReApplys_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 97:20]
  assign Broadcaster_io_remote_in_valid = ReScatter_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 93:28]
  assign Broadcaster_io_remote_in_bits_tdata = ReScatter_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 93:28]
  assign Broadcaster_io_remote_in_bits_tkeep = ReScatter_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 93:28]
  assign Broadcaster_io_local_fpga_id = controls_io_data_16[1:0]; // @[nf_arm_doce_top_main.scala 171:32]
  assign Broadcaster_io_flush = Scatters_0_io_issue_sync & Scatters_1_io_issue_sync & Scatters_2_io_issue_sync &
    Scatters_3_io_issue_sync; // @[nf_arm_doce_top_main.scala 172:70]
  assign Broadcaster_io_signal = controls_io_signal & controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 173:47]
  assign ReApplys_0_clock = clock;
  assign ReApplys_0_reset = reset;
  assign ReApplys_0_io_xbar_in_valid = Broadcaster_io_remote_out_0_valid; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_0_io_xbar_in_bits_tdata = Broadcaster_io_remote_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_0_io_xbar_in_bits_tkeep = Broadcaster_io_remote_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_0_io_remote_out_ready = ReSwitch_io_xbar_in_0_ready; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReApplys_0_io_recv_sync = {Scatters_0_io_recv_sync_hi_hi,ReApplys_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 150:75]
  assign ReApplys_0_io_recv_sync_phase2 = ReScatter_io_issue_sync_phase2_0; // @[nf_arm_doce_top_main.scala 154:29]
  assign ReApplys_0_io_signal = controls_io_signal & controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 152:41]
  assign ReApplys_0_io_local_fpga_id = controls_io_data_16[1:0]; // @[nf_arm_doce_top_main.scala 151:26]
  assign ReApplys_0_io_packet_size = controls_io_data_25; // @[nf_arm_doce_top_main.scala 155:24]
  assign ReApplys_0_io_level = controls_io_level; // @[nf_arm_doce_top_main.scala 156:18]
  assign ReApplys_0_io_pending_time = {{16'd0}, controls_io_data_26[15:0]}; // @[nf_arm_doce_top_main.scala 157:65]
  assign ReApplys_0_io_pending_parameter = {{16'd0}, controls_io_data_26[31:16]}; // @[nf_arm_doce_top_main.scala 158:70]
  assign ReApplys_0_io_idol_fpga_num = ReScatter_io_idol_fpga_num; // @[nf_arm_doce_top_main.scala 159:26]
  assign ReApplys_1_clock = clock;
  assign ReApplys_1_reset = reset;
  assign ReApplys_1_io_xbar_in_valid = Broadcaster_io_remote_out_1_valid; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_1_io_xbar_in_bits_tdata = Broadcaster_io_remote_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_1_io_xbar_in_bits_tkeep = Broadcaster_io_remote_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_1_io_remote_out_ready = ReSwitch_io_xbar_in_1_ready; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReApplys_1_io_recv_sync = {Scatters_0_io_recv_sync_hi_hi,ReApplys_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 150:75]
  assign ReApplys_1_io_recv_sync_phase2 = ReScatter_io_issue_sync_phase2_1; // @[nf_arm_doce_top_main.scala 154:29]
  assign ReApplys_1_io_signal = controls_io_signal & controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 152:41]
  assign ReApplys_1_io_local_fpga_id = controls_io_data_16[1:0]; // @[nf_arm_doce_top_main.scala 151:26]
  assign ReApplys_1_io_packet_size = controls_io_data_25; // @[nf_arm_doce_top_main.scala 155:24]
  assign ReApplys_1_io_level = controls_io_level; // @[nf_arm_doce_top_main.scala 156:18]
  assign ReApplys_1_io_pending_time = {{16'd0}, controls_io_data_26[15:0]}; // @[nf_arm_doce_top_main.scala 157:65]
  assign ReApplys_1_io_pending_parameter = {{16'd0}, controls_io_data_26[31:16]}; // @[nf_arm_doce_top_main.scala 158:70]
  assign ReApplys_1_io_idol_fpga_num = ReScatter_io_idol_fpga_num; // @[nf_arm_doce_top_main.scala 159:26]
  assign ReApplys_2_clock = clock;
  assign ReApplys_2_reset = reset;
  assign ReApplys_2_io_xbar_in_valid = Broadcaster_io_remote_out_2_valid; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_2_io_xbar_in_bits_tdata = Broadcaster_io_remote_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_2_io_xbar_in_bits_tkeep = Broadcaster_io_remote_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_2_io_remote_out_ready = ReSwitch_io_xbar_in_2_ready; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReApplys_2_io_recv_sync = {Scatters_0_io_recv_sync_hi_hi,ReApplys_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 150:75]
  assign ReApplys_2_io_recv_sync_phase2 = ReScatter_io_issue_sync_phase2_2; // @[nf_arm_doce_top_main.scala 154:29]
  assign ReApplys_2_io_signal = controls_io_signal & controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 152:41]
  assign ReApplys_2_io_local_fpga_id = controls_io_data_16[1:0]; // @[nf_arm_doce_top_main.scala 151:26]
  assign ReApplys_2_io_packet_size = controls_io_data_25; // @[nf_arm_doce_top_main.scala 155:24]
  assign ReApplys_2_io_level = controls_io_level; // @[nf_arm_doce_top_main.scala 156:18]
  assign ReApplys_2_io_pending_time = {{16'd0}, controls_io_data_26[15:0]}; // @[nf_arm_doce_top_main.scala 157:65]
  assign ReApplys_2_io_pending_parameter = {{16'd0}, controls_io_data_26[31:16]}; // @[nf_arm_doce_top_main.scala 158:70]
  assign ReApplys_2_io_idol_fpga_num = ReScatter_io_idol_fpga_num; // @[nf_arm_doce_top_main.scala 159:26]
  assign ReApplys_3_clock = clock;
  assign ReApplys_3_reset = reset;
  assign ReApplys_3_io_xbar_in_valid = Broadcaster_io_remote_out_3_valid; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_3_io_xbar_in_bits_tdata = Broadcaster_io_remote_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_3_io_xbar_in_bits_tkeep = Broadcaster_io_remote_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 97:20]
  assign ReApplys_3_io_remote_out_ready = ReSwitch_io_xbar_in_3_ready; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReApplys_3_io_recv_sync = {Scatters_0_io_recv_sync_hi_hi,ReApplys_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 150:75]
  assign ReApplys_3_io_recv_sync_phase2 = ReScatter_io_issue_sync_phase2_3; // @[nf_arm_doce_top_main.scala 154:29]
  assign ReApplys_3_io_signal = controls_io_signal & controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 152:41]
  assign ReApplys_3_io_local_fpga_id = controls_io_data_16[1:0]; // @[nf_arm_doce_top_main.scala 151:26]
  assign ReApplys_3_io_packet_size = controls_io_data_25; // @[nf_arm_doce_top_main.scala 155:24]
  assign ReApplys_3_io_level = controls_io_level; // @[nf_arm_doce_top_main.scala 156:18]
  assign ReApplys_3_io_pending_time = {{16'd0}, controls_io_data_26[15:0]}; // @[nf_arm_doce_top_main.scala 157:65]
  assign ReApplys_3_io_pending_parameter = {{16'd0}, controls_io_data_26[31:16]}; // @[nf_arm_doce_top_main.scala 158:70]
  assign ReApplys_3_io_idol_fpga_num = ReScatter_io_idol_fpga_num; // @[nf_arm_doce_top_main.scala 159:26]
  assign ReScatter_clock = clock;
  assign ReScatter_reset = reset;
  assign ReScatter_io_remote_in_w_valid = io_Re_memory_in_w_valid; // @[nf_arm_doce_top_main.scala 94:26]
  assign ReScatter_io_remote_in_w_bits_wdata = io_Re_memory_in_w_bits_wdata; // @[nf_arm_doce_top_main.scala 94:26]
  assign ReScatter_io_remote_in_w_bits_wstrb = io_Re_memory_in_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 94:26]
  assign ReScatter_io_xbar_out_ready = Broadcaster_io_remote_in_ready; // @[nf_arm_doce_top_main.scala 93:28]
  assign ReScatter_io_signal = controls_io_signal & controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 164:45]
  assign ReScatter_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 163:22]
  assign ReScatter_io_local_fpga_id = controls_io_data_16[1:0]; // @[nf_arm_doce_top_main.scala 165:30]
  assign ReSwitch_clock = clock;
  assign ReSwitch_reset = reset;
  assign ReSwitch_io_xbar_in_0_valid = ReApplys_0_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_0_bits_tdata = ReApplys_0_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_0_bits_tkeep = ReApplys_0_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_0_bits_tlast = ReApplys_0_io_remote_out_bits_tlast; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_1_valid = ReApplys_1_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_1_bits_tdata = ReApplys_1_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_1_bits_tkeep = ReApplys_1_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_1_bits_tlast = ReApplys_1_io_remote_out_bits_tlast; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_2_valid = ReApplys_2_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_2_bits_tdata = ReApplys_2_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_2_bits_tkeep = ReApplys_2_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_2_bits_tlast = ReApplys_2_io_remote_out_bits_tlast; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_3_valid = ReApplys_3_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_3_bits_tdata = ReApplys_3_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_3_bits_tkeep = ReApplys_3_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_xbar_in_3_bits_tlast = ReApplys_3_io_remote_out_bits_tlast; // @[nf_arm_doce_top_main.scala 98:30]
  assign ReSwitch_io_remote_out_aw_ready = io_Re_memory_out_aw_ready; // @[nf_arm_doce_top_main.scala 101:20]
  assign ReSwitch_io_remote_out_w_ready = io_Re_memory_out_w_ready; // @[nf_arm_doce_top_main.scala 101:20]
  assign ReSwitch_io_level_base_addr_0 = {controls_io_data_18,controls_io_data_17}; // @[Cat.scala 30:58]
  assign ReSwitch_io_level_base_addr_1 = {controls_io_data_20,controls_io_data_19}; // @[Cat.scala 30:58]
  assign ReSwitch_io_level_base_addr_2 = {controls_io_data_22,controls_io_data_21}; // @[Cat.scala 30:58]
  assign ReSwitch_io_level_base_addr_3 = {controls_io_data_24,controls_io_data_23}; // @[Cat.scala 30:58]
  assign ReSwitch_io_net_constrain = controls_io_data_27; // @[nf_arm_doce_top_main.scala 170:29]
  always @(posedge clock) begin
    if (reset) begin // @[nf_arm_doce_top_main.scala 59:32]
      max_size_to_net <= 32'h0; // @[nf_arm_doce_top_main.scala 59:32]
    end else if (!(io_Re_memory_out_w_valid & io_Re_memory_out_w_ready)) begin // @[nf_arm_doce_top_main.scala 62:79]
      if (controls_io_signal) begin // @[nf_arm_doce_top_main.scala 64:33]
        if (size_to_net > max_size_to_net) begin // @[nf_arm_doce_top_main.scala 66:40]
          max_size_to_net <= size_to_net; // @[nf_arm_doce_top_main.scala 67:23]
        end
      end
    end
    if (reset) begin // @[nf_arm_doce_top_main.scala 61:28]
      size_to_net <= 32'h0; // @[nf_arm_doce_top_main.scala 61:28]
    end else if (io_Re_memory_out_w_valid & io_Re_memory_out_w_ready) begin // @[nf_arm_doce_top_main.scala 62:79]
      size_to_net <= _size_to_net_T_1; // @[nf_arm_doce_top_main.scala 63:17]
    end else if (controls_io_signal) begin // @[nf_arm_doce_top_main.scala 64:33]
      size_to_net <= 32'h0; // @[nf_arm_doce_top_main.scala 65:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  max_size_to_net = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  size_to_net = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
