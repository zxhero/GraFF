module LookupTable(
  input         clock,
  input         reset,
  output [31:0] io_data_0,
  output [31:0] io_data_1,
  output [31:0] io_data_2,
  output [31:0] io_data_3,
  output [31:0] io_data_4,
  output [31:0] io_data_5,
  output [31:0] io_data_6,
  output [31:0] io_data_7,
  output [31:0] io_data_8,
  output [31:0] io_data_9,
  output [31:0] io_data_10,
  output [31:0] io_data_11,
  output [31:0] io_data_12,
  output [31:0] io_data_13,
  input  [31:0] io_dataIn_0,
  input  [31:0] io_dataIn_1,
  input         io_writeFlag_0,
  input         io_writeFlag_1,
  input  [4:0]  io_wptr_0,
  input  [4:0]  io_wptr_1,
  input  [63:0] config_awaddr,
  output        config_awready,
  input  [63:0] config_araddr,
  input         config_arvalid,
  output        config_arready,
  input  [31:0] config_wdata,
  input  [3:0]  config_wstrb,
  input         config_wvalid,
  output        config_wready,
  output [31:0] config_rdata,
  output        config_rvalid,
  input         config_rready,
  output        config_bvalid,
  input         config_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] table_0; // @[numa.scala 17:22]
  reg [31:0] table_1; // @[numa.scala 17:22]
  reg [31:0] table_2; // @[numa.scala 17:22]
  reg [31:0] table_3; // @[numa.scala 17:22]
  reg [31:0] table_4; // @[numa.scala 17:22]
  reg [31:0] table_5; // @[numa.scala 17:22]
  reg [31:0] table_6; // @[numa.scala 17:22]
  reg [31:0] table_7; // @[numa.scala 17:22]
  reg [31:0] table_8; // @[numa.scala 17:22]
  reg [31:0] table_9; // @[numa.scala 17:22]
  reg [31:0] table_10; // @[numa.scala 17:22]
  reg [31:0] table_11; // @[numa.scala 17:22]
  reg [31:0] table_12; // @[numa.scala 17:22]
  reg [31:0] table_13; // @[numa.scala 17:22]
  reg [31:0] table_14; // @[numa.scala 17:22]
  reg [31:0] table_15; // @[numa.scala 17:22]
  reg [31:0] table_16; // @[numa.scala 17:22]
  reg [31:0] table_17; // @[numa.scala 17:22]
  reg [31:0] table_18; // @[numa.scala 17:22]
  reg [31:0] table_19; // @[numa.scala 17:22]
  reg [31:0] table_20; // @[numa.scala 17:22]
  reg [31:0] table_21; // @[numa.scala 17:22]
  reg [31:0] table_22; // @[numa.scala 17:22]
  reg [31:0] table_23; // @[numa.scala 17:22]
  reg [31:0] table_24; // @[numa.scala 17:22]
  reg [31:0] table_25; // @[numa.scala 17:22]
  reg [31:0] table_26; // @[numa.scala 17:22]
  reg [31:0] table_27; // @[numa.scala 17:22]
  reg [31:0] table_28; // @[numa.scala 17:22]
  reg [31:0] table_29; // @[numa.scala 17:22]
  reg [31:0] table_30; // @[numa.scala 17:22]
  reg [31:0] table_31; // @[numa.scala 17:22]
  reg  rvalid; // @[numa.scala 18:23]
  reg  bvalid; // @[numa.scala 19:23]
  wire  _config_arready_T = ~rvalid; // @[numa.scala 25:28]
  wire [4:0] ewaddr = config_awaddr[6:2]; // @[numa.scala 65:26]
  wire [31:0] _GEN_1 = 5'h1 == ewaddr ? table_1 : table_0; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_2 = 5'h2 == ewaddr ? table_2 : _GEN_1; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_3 = 5'h3 == ewaddr ? table_3 : _GEN_2; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_4 = 5'h4 == ewaddr ? table_4 : _GEN_3; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_5 = 5'h5 == ewaddr ? table_5 : _GEN_4; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_6 = 5'h6 == ewaddr ? table_6 : _GEN_5; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_7 = 5'h7 == ewaddr ? table_7 : _GEN_6; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_8 = 5'h8 == ewaddr ? table_8 : _GEN_7; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_9 = 5'h9 == ewaddr ? table_9 : _GEN_8; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_10 = 5'ha == ewaddr ? table_10 : _GEN_9; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_11 = 5'hb == ewaddr ? table_11 : _GEN_10; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_12 = 5'hc == ewaddr ? table_12 : _GEN_11; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_13 = 5'hd == ewaddr ? table_13 : _GEN_12; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_14 = 5'he == ewaddr ? table_14 : _GEN_13; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_15 = 5'hf == ewaddr ? table_15 : _GEN_14; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_16 = 5'h10 == ewaddr ? table_16 : _GEN_15; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_17 = 5'h11 == ewaddr ? table_17 : _GEN_16; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_18 = 5'h12 == ewaddr ? table_18 : _GEN_17; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_19 = 5'h13 == ewaddr ? table_19 : _GEN_18; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_20 = 5'h14 == ewaddr ? table_20 : _GEN_19; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_21 = 5'h15 == ewaddr ? table_21 : _GEN_20; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_22 = 5'h16 == ewaddr ? table_22 : _GEN_21; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_23 = 5'h17 == ewaddr ? table_23 : _GEN_22; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_24 = 5'h18 == ewaddr ? table_24 : _GEN_23; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_25 = 5'h19 == ewaddr ? table_25 : _GEN_24; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_26 = 5'h1a == ewaddr ? table_26 : _GEN_25; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_27 = 5'h1b == ewaddr ? table_27 : _GEN_26; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_28 = 5'h1c == ewaddr ? table_28 : _GEN_27; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_29 = 5'h1d == ewaddr ? table_29 : _GEN_28; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_30 = 5'h1e == ewaddr ? table_30 : _GEN_29; // @[numa.scala 36:91 numa.scala 36:91]
  wire [31:0] _GEN_31 = 5'h1f == ewaddr ? table_31 : _GEN_30; // @[numa.scala 36:91 numa.scala 36:91]
  wire  wbytesvalid_0 = config_wvalid & config_wstrb[0]; // @[numa.scala 40:39]
  wire [7:0] wbytes_0 = wbytesvalid_0 ? config_wdata[7:0] : _GEN_31[7:0]; // @[numa.scala 36:29]
  wire  wbytesvalid_1 = config_wvalid & config_wstrb[1]; // @[numa.scala 40:39]
  wire [7:0] wbytes_1 = wbytesvalid_1 ? config_wdata[15:8] : _GEN_31[15:8]; // @[numa.scala 36:29]
  wire  wbytesvalid_2 = config_wvalid & config_wstrb[2]; // @[numa.scala 40:39]
  wire [7:0] wbytes_2 = wbytesvalid_2 ? config_wdata[23:16] : _GEN_31[23:16]; // @[numa.scala 36:29]
  wire  wbytesvalid_3 = config_wvalid & config_wstrb[3]; // @[numa.scala 40:39]
  wire [7:0] wbytes_3 = wbytesvalid_3 ? config_wdata[31:24] : _GEN_31[31:24]; // @[numa.scala 36:29]
  wire  _T = io_writeFlag_0 & io_writeFlag_1; // @[numa.scala 43:46]
  wire [31:0] _table_T = {wbytes_3,wbytes_2,wbytes_1,wbytes_0}; // @[numa.scala 44:35]
  wire [31:0] _GEN_32 = 5'h0 == ewaddr ? _table_T : table_0; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_33 = 5'h1 == ewaddr ? _table_T : table_1; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_34 = 5'h2 == ewaddr ? _table_T : table_2; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_35 = 5'h3 == ewaddr ? _table_T : table_3; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_36 = 5'h4 == ewaddr ? _table_T : table_4; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_37 = 5'h5 == ewaddr ? _table_T : table_5; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_38 = 5'h6 == ewaddr ? _table_T : table_6; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_39 = 5'h7 == ewaddr ? _table_T : table_7; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_40 = 5'h8 == ewaddr ? _table_T : table_8; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_41 = 5'h9 == ewaddr ? _table_T : table_9; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_42 = 5'ha == ewaddr ? _table_T : table_10; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_43 = 5'hb == ewaddr ? _table_T : table_11; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_44 = 5'hc == ewaddr ? _table_T : table_12; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_45 = 5'hd == ewaddr ? _table_T : table_13; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_46 = 5'he == ewaddr ? _table_T : table_14; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_47 = 5'hf == ewaddr ? _table_T : table_15; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_48 = 5'h10 == ewaddr ? _table_T : table_16; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_49 = 5'h11 == ewaddr ? _table_T : table_17; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_50 = 5'h12 == ewaddr ? _table_T : table_18; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_51 = 5'h13 == ewaddr ? _table_T : table_19; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_52 = 5'h14 == ewaddr ? _table_T : table_20; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_53 = 5'h15 == ewaddr ? _table_T : table_21; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_54 = 5'h16 == ewaddr ? _table_T : table_22; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_55 = 5'h17 == ewaddr ? _table_T : table_23; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_56 = 5'h18 == ewaddr ? _table_T : table_24; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_57 = 5'h19 == ewaddr ? _table_T : table_25; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_58 = 5'h1a == ewaddr ? _table_T : table_26; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_59 = 5'h1b == ewaddr ? _table_T : table_27; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_60 = 5'h1c == ewaddr ? _table_T : table_28; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_61 = 5'h1d == ewaddr ? _table_T : table_29; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_62 = 5'h1e == ewaddr ? _table_T : table_30; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_63 = 5'h1f == ewaddr ? _table_T : table_31; // @[numa.scala 44:19 numa.scala 44:19 numa.scala 17:22]
  wire [31:0] _GEN_64 = 5'h0 == io_wptr_0 ? io_dataIn_0 : _GEN_32; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_65 = 5'h1 == io_wptr_0 ? io_dataIn_0 : _GEN_33; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_66 = 5'h2 == io_wptr_0 ? io_dataIn_0 : _GEN_34; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_67 = 5'h3 == io_wptr_0 ? io_dataIn_0 : _GEN_35; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_68 = 5'h4 == io_wptr_0 ? io_dataIn_0 : _GEN_36; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_69 = 5'h5 == io_wptr_0 ? io_dataIn_0 : _GEN_37; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_70 = 5'h6 == io_wptr_0 ? io_dataIn_0 : _GEN_38; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_71 = 5'h7 == io_wptr_0 ? io_dataIn_0 : _GEN_39; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_72 = 5'h8 == io_wptr_0 ? io_dataIn_0 : _GEN_40; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_73 = 5'h9 == io_wptr_0 ? io_dataIn_0 : _GEN_41; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_74 = 5'ha == io_wptr_0 ? io_dataIn_0 : _GEN_42; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_75 = 5'hb == io_wptr_0 ? io_dataIn_0 : _GEN_43; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_76 = 5'hc == io_wptr_0 ? io_dataIn_0 : _GEN_44; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_77 = 5'hd == io_wptr_0 ? io_dataIn_0 : _GEN_45; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_78 = 5'he == io_wptr_0 ? io_dataIn_0 : _GEN_46; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_79 = 5'hf == io_wptr_0 ? io_dataIn_0 : _GEN_47; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_80 = 5'h10 == io_wptr_0 ? io_dataIn_0 : _GEN_48; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_81 = 5'h11 == io_wptr_0 ? io_dataIn_0 : _GEN_49; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_82 = 5'h12 == io_wptr_0 ? io_dataIn_0 : _GEN_50; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_83 = 5'h13 == io_wptr_0 ? io_dataIn_0 : _GEN_51; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_84 = 5'h14 == io_wptr_0 ? io_dataIn_0 : _GEN_52; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_85 = 5'h15 == io_wptr_0 ? io_dataIn_0 : _GEN_53; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_86 = 5'h16 == io_wptr_0 ? io_dataIn_0 : _GEN_54; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_87 = 5'h17 == io_wptr_0 ? io_dataIn_0 : _GEN_55; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_88 = 5'h18 == io_wptr_0 ? io_dataIn_0 : _GEN_56; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_89 = 5'h19 == io_wptr_0 ? io_dataIn_0 : _GEN_57; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_90 = 5'h1a == io_wptr_0 ? io_dataIn_0 : _GEN_58; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_91 = 5'h1b == io_wptr_0 ? io_dataIn_0 : _GEN_59; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_92 = 5'h1c == io_wptr_0 ? io_dataIn_0 : _GEN_60; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_93 = 5'h1d == io_wptr_0 ? io_dataIn_0 : _GEN_61; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_94 = 5'h1e == io_wptr_0 ? io_dataIn_0 : _GEN_62; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_95 = 5'h1f == io_wptr_0 ? io_dataIn_0 : _GEN_63; // @[numa.scala 45:23 numa.scala 45:23]
  wire [31:0] _GEN_224 = 5'h0 == io_wptr_1 ? io_dataIn_1 : _GEN_32; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_225 = 5'h1 == io_wptr_1 ? io_dataIn_1 : _GEN_33; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_226 = 5'h2 == io_wptr_1 ? io_dataIn_1 : _GEN_34; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_227 = 5'h3 == io_wptr_1 ? io_dataIn_1 : _GEN_35; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_228 = 5'h4 == io_wptr_1 ? io_dataIn_1 : _GEN_36; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_229 = 5'h5 == io_wptr_1 ? io_dataIn_1 : _GEN_37; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_230 = 5'h6 == io_wptr_1 ? io_dataIn_1 : _GEN_38; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_231 = 5'h7 == io_wptr_1 ? io_dataIn_1 : _GEN_39; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_232 = 5'h8 == io_wptr_1 ? io_dataIn_1 : _GEN_40; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_233 = 5'h9 == io_wptr_1 ? io_dataIn_1 : _GEN_41; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_234 = 5'ha == io_wptr_1 ? io_dataIn_1 : _GEN_42; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_235 = 5'hb == io_wptr_1 ? io_dataIn_1 : _GEN_43; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_236 = 5'hc == io_wptr_1 ? io_dataIn_1 : _GEN_44; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_237 = 5'hd == io_wptr_1 ? io_dataIn_1 : _GEN_45; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_238 = 5'he == io_wptr_1 ? io_dataIn_1 : _GEN_46; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_239 = 5'hf == io_wptr_1 ? io_dataIn_1 : _GEN_47; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_240 = 5'h10 == io_wptr_1 ? io_dataIn_1 : _GEN_48; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_241 = 5'h11 == io_wptr_1 ? io_dataIn_1 : _GEN_49; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_242 = 5'h12 == io_wptr_1 ? io_dataIn_1 : _GEN_50; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_243 = 5'h13 == io_wptr_1 ? io_dataIn_1 : _GEN_51; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_244 = 5'h14 == io_wptr_1 ? io_dataIn_1 : _GEN_52; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_245 = 5'h15 == io_wptr_1 ? io_dataIn_1 : _GEN_53; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_246 = 5'h16 == io_wptr_1 ? io_dataIn_1 : _GEN_54; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_247 = 5'h17 == io_wptr_1 ? io_dataIn_1 : _GEN_55; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_248 = 5'h18 == io_wptr_1 ? io_dataIn_1 : _GEN_56; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_249 = 5'h19 == io_wptr_1 ? io_dataIn_1 : _GEN_57; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_250 = 5'h1a == io_wptr_1 ? io_dataIn_1 : _GEN_58; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_251 = 5'h1b == io_wptr_1 ? io_dataIn_1 : _GEN_59; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_252 = 5'h1c == io_wptr_1 ? io_dataIn_1 : _GEN_60; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_253 = 5'h1d == io_wptr_1 ? io_dataIn_1 : _GEN_61; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_254 = 5'h1e == io_wptr_1 ? io_dataIn_1 : _GEN_62; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_255 = 5'h1f == io_wptr_1 ? io_dataIn_1 : _GEN_63; // @[numa.scala 52:23 numa.scala 52:23]
  wire [31:0] _GEN_288 = 5'h0 == io_wptr_0 ? io_dataIn_0 : table_0; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_289 = 5'h1 == io_wptr_0 ? io_dataIn_0 : table_1; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_290 = 5'h2 == io_wptr_0 ? io_dataIn_0 : table_2; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_291 = 5'h3 == io_wptr_0 ? io_dataIn_0 : table_3; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_292 = 5'h4 == io_wptr_0 ? io_dataIn_0 : table_4; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_293 = 5'h5 == io_wptr_0 ? io_dataIn_0 : table_5; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_294 = 5'h6 == io_wptr_0 ? io_dataIn_0 : table_6; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_295 = 5'h7 == io_wptr_0 ? io_dataIn_0 : table_7; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_296 = 5'h8 == io_wptr_0 ? io_dataIn_0 : table_8; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_297 = 5'h9 == io_wptr_0 ? io_dataIn_0 : table_9; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_298 = 5'ha == io_wptr_0 ? io_dataIn_0 : table_10; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_299 = 5'hb == io_wptr_0 ? io_dataIn_0 : table_11; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_300 = 5'hc == io_wptr_0 ? io_dataIn_0 : table_12; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_301 = 5'hd == io_wptr_0 ? io_dataIn_0 : table_13; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_302 = 5'he == io_wptr_0 ? io_dataIn_0 : table_14; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_303 = 5'hf == io_wptr_0 ? io_dataIn_0 : table_15; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_304 = 5'h10 == io_wptr_0 ? io_dataIn_0 : table_16; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_305 = 5'h11 == io_wptr_0 ? io_dataIn_0 : table_17; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_306 = 5'h12 == io_wptr_0 ? io_dataIn_0 : table_18; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_307 = 5'h13 == io_wptr_0 ? io_dataIn_0 : table_19; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_308 = 5'h14 == io_wptr_0 ? io_dataIn_0 : table_20; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_309 = 5'h15 == io_wptr_0 ? io_dataIn_0 : table_21; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_310 = 5'h16 == io_wptr_0 ? io_dataIn_0 : table_22; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_311 = 5'h17 == io_wptr_0 ? io_dataIn_0 : table_23; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_312 = 5'h18 == io_wptr_0 ? io_dataIn_0 : table_24; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_313 = 5'h19 == io_wptr_0 ? io_dataIn_0 : table_25; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_314 = 5'h1a == io_wptr_0 ? io_dataIn_0 : table_26; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_315 = 5'h1b == io_wptr_0 ? io_dataIn_0 : table_27; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_316 = 5'h1c == io_wptr_0 ? io_dataIn_0 : table_28; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_317 = 5'h1d == io_wptr_0 ? io_dataIn_0 : table_29; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_318 = 5'h1e == io_wptr_0 ? io_dataIn_0 : table_30; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_319 = 5'h1f == io_wptr_0 ? io_dataIn_0 : table_31; // @[numa.scala 56:23 numa.scala 56:23 numa.scala 17:22]
  wire [31:0] _GEN_320 = 5'h0 == io_wptr_1 ? io_dataIn_1 : _GEN_288; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_321 = 5'h1 == io_wptr_1 ? io_dataIn_1 : _GEN_289; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_322 = 5'h2 == io_wptr_1 ? io_dataIn_1 : _GEN_290; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_323 = 5'h3 == io_wptr_1 ? io_dataIn_1 : _GEN_291; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_324 = 5'h4 == io_wptr_1 ? io_dataIn_1 : _GEN_292; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_325 = 5'h5 == io_wptr_1 ? io_dataIn_1 : _GEN_293; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_326 = 5'h6 == io_wptr_1 ? io_dataIn_1 : _GEN_294; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_327 = 5'h7 == io_wptr_1 ? io_dataIn_1 : _GEN_295; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_328 = 5'h8 == io_wptr_1 ? io_dataIn_1 : _GEN_296; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_329 = 5'h9 == io_wptr_1 ? io_dataIn_1 : _GEN_297; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_330 = 5'ha == io_wptr_1 ? io_dataIn_1 : _GEN_298; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_331 = 5'hb == io_wptr_1 ? io_dataIn_1 : _GEN_299; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_332 = 5'hc == io_wptr_1 ? io_dataIn_1 : _GEN_300; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_333 = 5'hd == io_wptr_1 ? io_dataIn_1 : _GEN_301; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_334 = 5'he == io_wptr_1 ? io_dataIn_1 : _GEN_302; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_335 = 5'hf == io_wptr_1 ? io_dataIn_1 : _GEN_303; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_336 = 5'h10 == io_wptr_1 ? io_dataIn_1 : _GEN_304; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_337 = 5'h11 == io_wptr_1 ? io_dataIn_1 : _GEN_305; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_338 = 5'h12 == io_wptr_1 ? io_dataIn_1 : _GEN_306; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_339 = 5'h13 == io_wptr_1 ? io_dataIn_1 : _GEN_307; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_340 = 5'h14 == io_wptr_1 ? io_dataIn_1 : _GEN_308; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_341 = 5'h15 == io_wptr_1 ? io_dataIn_1 : _GEN_309; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_342 = 5'h16 == io_wptr_1 ? io_dataIn_1 : _GEN_310; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_343 = 5'h17 == io_wptr_1 ? io_dataIn_1 : _GEN_311; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_344 = 5'h18 == io_wptr_1 ? io_dataIn_1 : _GEN_312; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_345 = 5'h19 == io_wptr_1 ? io_dataIn_1 : _GEN_313; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_346 = 5'h1a == io_wptr_1 ? io_dataIn_1 : _GEN_314; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_347 = 5'h1b == io_wptr_1 ? io_dataIn_1 : _GEN_315; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_348 = 5'h1c == io_wptr_1 ? io_dataIn_1 : _GEN_316; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_349 = 5'h1d == io_wptr_1 ? io_dataIn_1 : _GEN_317; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_350 = 5'h1e == io_wptr_1 ? io_dataIn_1 : _GEN_318; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_351 = 5'h1f == io_wptr_1 ? io_dataIn_1 : _GEN_319; // @[numa.scala 57:23 numa.scala 57:23]
  wire [31:0] _GEN_384 = 5'h0 == io_wptr_1 ? io_dataIn_1 : table_0; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_385 = 5'h1 == io_wptr_1 ? io_dataIn_1 : table_1; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_386 = 5'h2 == io_wptr_1 ? io_dataIn_1 : table_2; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_387 = 5'h3 == io_wptr_1 ? io_dataIn_1 : table_3; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_388 = 5'h4 == io_wptr_1 ? io_dataIn_1 : table_4; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_389 = 5'h5 == io_wptr_1 ? io_dataIn_1 : table_5; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_390 = 5'h6 == io_wptr_1 ? io_dataIn_1 : table_6; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_391 = 5'h7 == io_wptr_1 ? io_dataIn_1 : table_7; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_392 = 5'h8 == io_wptr_1 ? io_dataIn_1 : table_8; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_393 = 5'h9 == io_wptr_1 ? io_dataIn_1 : table_9; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_394 = 5'ha == io_wptr_1 ? io_dataIn_1 : table_10; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_395 = 5'hb == io_wptr_1 ? io_dataIn_1 : table_11; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_396 = 5'hc == io_wptr_1 ? io_dataIn_1 : table_12; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_397 = 5'hd == io_wptr_1 ? io_dataIn_1 : table_13; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_398 = 5'he == io_wptr_1 ? io_dataIn_1 : table_14; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_399 = 5'hf == io_wptr_1 ? io_dataIn_1 : table_15; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_400 = 5'h10 == io_wptr_1 ? io_dataIn_1 : table_16; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_401 = 5'h11 == io_wptr_1 ? io_dataIn_1 : table_17; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_402 = 5'h12 == io_wptr_1 ? io_dataIn_1 : table_18; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_403 = 5'h13 == io_wptr_1 ? io_dataIn_1 : table_19; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_404 = 5'h14 == io_wptr_1 ? io_dataIn_1 : table_20; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_405 = 5'h15 == io_wptr_1 ? io_dataIn_1 : table_21; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_406 = 5'h16 == io_wptr_1 ? io_dataIn_1 : table_22; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_407 = 5'h17 == io_wptr_1 ? io_dataIn_1 : table_23; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_408 = 5'h18 == io_wptr_1 ? io_dataIn_1 : table_24; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_409 = 5'h19 == io_wptr_1 ? io_dataIn_1 : table_25; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_410 = 5'h1a == io_wptr_1 ? io_dataIn_1 : table_26; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_411 = 5'h1b == io_wptr_1 ? io_dataIn_1 : table_27; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_412 = 5'h1c == io_wptr_1 ? io_dataIn_1 : table_28; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_413 = 5'h1d == io_wptr_1 ? io_dataIn_1 : table_29; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_414 = 5'h1e == io_wptr_1 ? io_dataIn_1 : table_30; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_415 = 5'h1f == io_wptr_1 ? io_dataIn_1 : table_31; // @[numa.scala 61:23 numa.scala 61:23 numa.scala 17:22]
  wire [31:0] _GEN_416 = io_writeFlag_1 ? _GEN_384 : table_0; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_417 = io_writeFlag_1 ? _GEN_385 : table_1; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_418 = io_writeFlag_1 ? _GEN_386 : table_2; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_419 = io_writeFlag_1 ? _GEN_387 : table_3; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_420 = io_writeFlag_1 ? _GEN_388 : table_4; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_421 = io_writeFlag_1 ? _GEN_389 : table_5; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_422 = io_writeFlag_1 ? _GEN_390 : table_6; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_423 = io_writeFlag_1 ? _GEN_391 : table_7; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_424 = io_writeFlag_1 ? _GEN_392 : table_8; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_425 = io_writeFlag_1 ? _GEN_393 : table_9; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_426 = io_writeFlag_1 ? _GEN_394 : table_10; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_427 = io_writeFlag_1 ? _GEN_395 : table_11; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_428 = io_writeFlag_1 ? _GEN_396 : table_12; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_429 = io_writeFlag_1 ? _GEN_397 : table_13; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_430 = io_writeFlag_1 ? _GEN_398 : table_14; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_431 = io_writeFlag_1 ? _GEN_399 : table_15; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_432 = io_writeFlag_1 ? _GEN_400 : table_16; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_433 = io_writeFlag_1 ? _GEN_401 : table_17; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_434 = io_writeFlag_1 ? _GEN_402 : table_18; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_435 = io_writeFlag_1 ? _GEN_403 : table_19; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_436 = io_writeFlag_1 ? _GEN_404 : table_20; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_437 = io_writeFlag_1 ? _GEN_405 : table_21; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_438 = io_writeFlag_1 ? _GEN_406 : table_22; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_439 = io_writeFlag_1 ? _GEN_407 : table_23; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_440 = io_writeFlag_1 ? _GEN_408 : table_24; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_441 = io_writeFlag_1 ? _GEN_409 : table_25; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_442 = io_writeFlag_1 ? _GEN_410 : table_26; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_443 = io_writeFlag_1 ? _GEN_411 : table_27; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_444 = io_writeFlag_1 ? _GEN_412 : table_28; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_445 = io_writeFlag_1 ? _GEN_413 : table_29; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_446 = io_writeFlag_1 ? _GEN_414 : table_30; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_447 = io_writeFlag_1 ? _GEN_415 : table_31; // @[numa.scala 60:30 numa.scala 17:22]
  wire [31:0] _GEN_448 = io_writeFlag_0 ? _GEN_288 : _GEN_416; // @[numa.scala 58:30]
  wire [31:0] _GEN_449 = io_writeFlag_0 ? _GEN_289 : _GEN_417; // @[numa.scala 58:30]
  wire [31:0] _GEN_450 = io_writeFlag_0 ? _GEN_290 : _GEN_418; // @[numa.scala 58:30]
  wire [31:0] _GEN_451 = io_writeFlag_0 ? _GEN_291 : _GEN_419; // @[numa.scala 58:30]
  wire [31:0] _GEN_452 = io_writeFlag_0 ? _GEN_292 : _GEN_420; // @[numa.scala 58:30]
  wire [31:0] _GEN_453 = io_writeFlag_0 ? _GEN_293 : _GEN_421; // @[numa.scala 58:30]
  wire [31:0] _GEN_454 = io_writeFlag_0 ? _GEN_294 : _GEN_422; // @[numa.scala 58:30]
  wire [31:0] _GEN_455 = io_writeFlag_0 ? _GEN_295 : _GEN_423; // @[numa.scala 58:30]
  wire [31:0] _GEN_456 = io_writeFlag_0 ? _GEN_296 : _GEN_424; // @[numa.scala 58:30]
  wire [31:0] _GEN_457 = io_writeFlag_0 ? _GEN_297 : _GEN_425; // @[numa.scala 58:30]
  wire [31:0] _GEN_458 = io_writeFlag_0 ? _GEN_298 : _GEN_426; // @[numa.scala 58:30]
  wire [31:0] _GEN_459 = io_writeFlag_0 ? _GEN_299 : _GEN_427; // @[numa.scala 58:30]
  wire [31:0] _GEN_460 = io_writeFlag_0 ? _GEN_300 : _GEN_428; // @[numa.scala 58:30]
  wire [31:0] _GEN_461 = io_writeFlag_0 ? _GEN_301 : _GEN_429; // @[numa.scala 58:30]
  wire [31:0] _GEN_462 = io_writeFlag_0 ? _GEN_302 : _GEN_430; // @[numa.scala 58:30]
  wire [31:0] _GEN_463 = io_writeFlag_0 ? _GEN_303 : _GEN_431; // @[numa.scala 58:30]
  wire [31:0] _GEN_464 = io_writeFlag_0 ? _GEN_304 : _GEN_432; // @[numa.scala 58:30]
  wire [31:0] _GEN_465 = io_writeFlag_0 ? _GEN_305 : _GEN_433; // @[numa.scala 58:30]
  wire [31:0] _GEN_466 = io_writeFlag_0 ? _GEN_306 : _GEN_434; // @[numa.scala 58:30]
  wire [31:0] _GEN_467 = io_writeFlag_0 ? _GEN_307 : _GEN_435; // @[numa.scala 58:30]
  wire [31:0] _GEN_468 = io_writeFlag_0 ? _GEN_308 : _GEN_436; // @[numa.scala 58:30]
  wire [31:0] _GEN_469 = io_writeFlag_0 ? _GEN_309 : _GEN_437; // @[numa.scala 58:30]
  wire [31:0] _GEN_470 = io_writeFlag_0 ? _GEN_310 : _GEN_438; // @[numa.scala 58:30]
  wire [31:0] _GEN_471 = io_writeFlag_0 ? _GEN_311 : _GEN_439; // @[numa.scala 58:30]
  wire [31:0] _GEN_472 = io_writeFlag_0 ? _GEN_312 : _GEN_440; // @[numa.scala 58:30]
  wire [31:0] _GEN_473 = io_writeFlag_0 ? _GEN_313 : _GEN_441; // @[numa.scala 58:30]
  wire [31:0] _GEN_474 = io_writeFlag_0 ? _GEN_314 : _GEN_442; // @[numa.scala 58:30]
  wire [31:0] _GEN_475 = io_writeFlag_0 ? _GEN_315 : _GEN_443; // @[numa.scala 58:30]
  wire [31:0] _GEN_476 = io_writeFlag_0 ? _GEN_316 : _GEN_444; // @[numa.scala 58:30]
  wire [31:0] _GEN_477 = io_writeFlag_0 ? _GEN_317 : _GEN_445; // @[numa.scala 58:30]
  wire [31:0] _GEN_478 = io_writeFlag_0 ? _GEN_318 : _GEN_446; // @[numa.scala 58:30]
  wire [31:0] _GEN_479 = io_writeFlag_0 ? _GEN_319 : _GEN_447; // @[numa.scala 58:30]
  wire [31:0] _GEN_480 = _T ? _GEN_320 : _GEN_448; // @[numa.scala 55:39]
  wire [31:0] _GEN_481 = _T ? _GEN_321 : _GEN_449; // @[numa.scala 55:39]
  wire [31:0] _GEN_482 = _T ? _GEN_322 : _GEN_450; // @[numa.scala 55:39]
  wire [31:0] _GEN_483 = _T ? _GEN_323 : _GEN_451; // @[numa.scala 55:39]
  wire [31:0] _GEN_484 = _T ? _GEN_324 : _GEN_452; // @[numa.scala 55:39]
  wire [31:0] _GEN_485 = _T ? _GEN_325 : _GEN_453; // @[numa.scala 55:39]
  wire [31:0] _GEN_486 = _T ? _GEN_326 : _GEN_454; // @[numa.scala 55:39]
  wire [31:0] _GEN_487 = _T ? _GEN_327 : _GEN_455; // @[numa.scala 55:39]
  wire [31:0] _GEN_488 = _T ? _GEN_328 : _GEN_456; // @[numa.scala 55:39]
  wire [31:0] _GEN_489 = _T ? _GEN_329 : _GEN_457; // @[numa.scala 55:39]
  wire [31:0] _GEN_490 = _T ? _GEN_330 : _GEN_458; // @[numa.scala 55:39]
  wire [31:0] _GEN_491 = _T ? _GEN_331 : _GEN_459; // @[numa.scala 55:39]
  wire [31:0] _GEN_492 = _T ? _GEN_332 : _GEN_460; // @[numa.scala 55:39]
  wire [31:0] _GEN_493 = _T ? _GEN_333 : _GEN_461; // @[numa.scala 55:39]
  wire [31:0] _GEN_494 = _T ? _GEN_334 : _GEN_462; // @[numa.scala 55:39]
  wire [31:0] _GEN_495 = _T ? _GEN_335 : _GEN_463; // @[numa.scala 55:39]
  wire [31:0] _GEN_496 = _T ? _GEN_336 : _GEN_464; // @[numa.scala 55:39]
  wire [31:0] _GEN_497 = _T ? _GEN_337 : _GEN_465; // @[numa.scala 55:39]
  wire [31:0] _GEN_498 = _T ? _GEN_338 : _GEN_466; // @[numa.scala 55:39]
  wire [31:0] _GEN_499 = _T ? _GEN_339 : _GEN_467; // @[numa.scala 55:39]
  wire [31:0] _GEN_500 = _T ? _GEN_340 : _GEN_468; // @[numa.scala 55:39]
  wire [31:0] _GEN_501 = _T ? _GEN_341 : _GEN_469; // @[numa.scala 55:39]
  wire [31:0] _GEN_502 = _T ? _GEN_342 : _GEN_470; // @[numa.scala 55:39]
  wire [31:0] _GEN_503 = _T ? _GEN_343 : _GEN_471; // @[numa.scala 55:39]
  wire [31:0] _GEN_504 = _T ? _GEN_344 : _GEN_472; // @[numa.scala 55:39]
  wire [31:0] _GEN_505 = _T ? _GEN_345 : _GEN_473; // @[numa.scala 55:39]
  wire [31:0] _GEN_506 = _T ? _GEN_346 : _GEN_474; // @[numa.scala 55:39]
  wire [31:0] _GEN_507 = _T ? _GEN_347 : _GEN_475; // @[numa.scala 55:39]
  wire [31:0] _GEN_508 = _T ? _GEN_348 : _GEN_476; // @[numa.scala 55:39]
  wire [31:0] _GEN_509 = _T ? _GEN_349 : _GEN_477; // @[numa.scala 55:39]
  wire [31:0] _GEN_510 = _T ? _GEN_350 : _GEN_478; // @[numa.scala 55:39]
  wire [31:0] _GEN_511 = _T ? _GEN_351 : _GEN_479; // @[numa.scala 55:39]
  wire [31:0] _GEN_512 = config_wvalid ? _GEN_32 : _GEN_480; // @[numa.scala 53:28]
  wire [31:0] _GEN_513 = config_wvalid ? _GEN_33 : _GEN_481; // @[numa.scala 53:28]
  wire [31:0] _GEN_514 = config_wvalid ? _GEN_34 : _GEN_482; // @[numa.scala 53:28]
  wire [31:0] _GEN_515 = config_wvalid ? _GEN_35 : _GEN_483; // @[numa.scala 53:28]
  wire [31:0] _GEN_516 = config_wvalid ? _GEN_36 : _GEN_484; // @[numa.scala 53:28]
  wire [31:0] _GEN_517 = config_wvalid ? _GEN_37 : _GEN_485; // @[numa.scala 53:28]
  wire [31:0] _GEN_518 = config_wvalid ? _GEN_38 : _GEN_486; // @[numa.scala 53:28]
  wire [31:0] _GEN_519 = config_wvalid ? _GEN_39 : _GEN_487; // @[numa.scala 53:28]
  wire [31:0] _GEN_520 = config_wvalid ? _GEN_40 : _GEN_488; // @[numa.scala 53:28]
  wire [31:0] _GEN_521 = config_wvalid ? _GEN_41 : _GEN_489; // @[numa.scala 53:28]
  wire [31:0] _GEN_522 = config_wvalid ? _GEN_42 : _GEN_490; // @[numa.scala 53:28]
  wire [31:0] _GEN_523 = config_wvalid ? _GEN_43 : _GEN_491; // @[numa.scala 53:28]
  wire [31:0] _GEN_524 = config_wvalid ? _GEN_44 : _GEN_492; // @[numa.scala 53:28]
  wire [31:0] _GEN_525 = config_wvalid ? _GEN_45 : _GEN_493; // @[numa.scala 53:28]
  wire [31:0] _GEN_526 = config_wvalid ? _GEN_46 : _GEN_494; // @[numa.scala 53:28]
  wire [31:0] _GEN_527 = config_wvalid ? _GEN_47 : _GEN_495; // @[numa.scala 53:28]
  wire [31:0] _GEN_528 = config_wvalid ? _GEN_48 : _GEN_496; // @[numa.scala 53:28]
  wire [31:0] _GEN_529 = config_wvalid ? _GEN_49 : _GEN_497; // @[numa.scala 53:28]
  wire [31:0] _GEN_530 = config_wvalid ? _GEN_50 : _GEN_498; // @[numa.scala 53:28]
  wire [31:0] _GEN_531 = config_wvalid ? _GEN_51 : _GEN_499; // @[numa.scala 53:28]
  wire [31:0] _GEN_532 = config_wvalid ? _GEN_52 : _GEN_500; // @[numa.scala 53:28]
  wire [31:0] _GEN_533 = config_wvalid ? _GEN_53 : _GEN_501; // @[numa.scala 53:28]
  wire [31:0] _GEN_534 = config_wvalid ? _GEN_54 : _GEN_502; // @[numa.scala 53:28]
  wire [31:0] _GEN_535 = config_wvalid ? _GEN_55 : _GEN_503; // @[numa.scala 53:28]
  wire [31:0] _GEN_536 = config_wvalid ? _GEN_56 : _GEN_504; // @[numa.scala 53:28]
  wire [31:0] _GEN_537 = config_wvalid ? _GEN_57 : _GEN_505; // @[numa.scala 53:28]
  wire [31:0] _GEN_538 = config_wvalid ? _GEN_58 : _GEN_506; // @[numa.scala 53:28]
  wire [31:0] _GEN_539 = config_wvalid ? _GEN_59 : _GEN_507; // @[numa.scala 53:28]
  wire [31:0] _GEN_540 = config_wvalid ? _GEN_60 : _GEN_508; // @[numa.scala 53:28]
  wire [31:0] _GEN_541 = config_wvalid ? _GEN_61 : _GEN_509; // @[numa.scala 53:28]
  wire [31:0] _GEN_542 = config_wvalid ? _GEN_62 : _GEN_510; // @[numa.scala 53:28]
  wire [31:0] _GEN_543 = config_wvalid ? _GEN_63 : _GEN_511; // @[numa.scala 53:28]
  reg [4:0] eraddr; // @[numa.scala 68:19]
  wire [31:0] _GEN_642 = 5'h1 == eraddr ? table_1 : table_0; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_643 = 5'h2 == eraddr ? table_2 : _GEN_642; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_644 = 5'h3 == eraddr ? table_3 : _GEN_643; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_645 = 5'h4 == eraddr ? table_4 : _GEN_644; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_646 = 5'h5 == eraddr ? table_5 : _GEN_645; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_647 = 5'h6 == eraddr ? table_6 : _GEN_646; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_648 = 5'h7 == eraddr ? table_7 : _GEN_647; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_649 = 5'h8 == eraddr ? table_8 : _GEN_648; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_650 = 5'h9 == eraddr ? table_9 : _GEN_649; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_651 = 5'ha == eraddr ? table_10 : _GEN_650; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_652 = 5'hb == eraddr ? table_11 : _GEN_651; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_653 = 5'hc == eraddr ? table_12 : _GEN_652; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_654 = 5'hd == eraddr ? table_13 : _GEN_653; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_655 = 5'he == eraddr ? table_14 : _GEN_654; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_656 = 5'hf == eraddr ? table_15 : _GEN_655; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_657 = 5'h10 == eraddr ? table_16 : _GEN_656; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_658 = 5'h11 == eraddr ? table_17 : _GEN_657; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_659 = 5'h12 == eraddr ? table_18 : _GEN_658; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_660 = 5'h13 == eraddr ? table_19 : _GEN_659; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_661 = 5'h14 == eraddr ? table_20 : _GEN_660; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_662 = 5'h15 == eraddr ? table_21 : _GEN_661; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_663 = 5'h16 == eraddr ? table_22 : _GEN_662; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_664 = 5'h17 == eraddr ? table_23 : _GEN_663; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_665 = 5'h18 == eraddr ? table_24 : _GEN_664; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_666 = 5'h19 == eraddr ? table_25 : _GEN_665; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_667 = 5'h1a == eraddr ? table_26 : _GEN_666; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_668 = 5'h1b == eraddr ? table_27 : _GEN_667; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_669 = 5'h1c == eraddr ? table_28 : _GEN_668; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_670 = 5'h1d == eraddr ? table_29 : _GEN_669; // @[numa.scala 76:16 numa.scala 76:16]
  wire [31:0] _GEN_671 = 5'h1e == eraddr ? table_30 : _GEN_670; // @[numa.scala 76:16 numa.scala 76:16]
  wire  _GEN_673 = rvalid & config_rready ? 1'h0 : rvalid; // @[numa.scala 80:38 numa.scala 81:12 numa.scala 18:23]
  wire  _GEN_674 = config_arvalid & _config_arready_T | _GEN_673; // @[numa.scala 78:45 numa.scala 79:12]
  wire  _GEN_675 = bvalid & config_bready ? 1'h0 : bvalid; // @[numa.scala 87:38 numa.scala 88:12 numa.scala 19:23]
  wire  _GEN_676 = config_wvalid | _GEN_675; // @[numa.scala 85:22 numa.scala 86:12]
  assign io_data_0 = table_0; // @[numa.scala 22:11]
  assign io_data_1 = table_1; // @[numa.scala 22:11]
  assign io_data_2 = table_2; // @[numa.scala 22:11]
  assign io_data_3 = table_3; // @[numa.scala 22:11]
  assign io_data_4 = table_4; // @[numa.scala 22:11]
  assign io_data_5 = table_5; // @[numa.scala 22:11]
  assign io_data_6 = table_6; // @[numa.scala 22:11]
  assign io_data_7 = table_7; // @[numa.scala 22:11]
  assign io_data_8 = table_8; // @[numa.scala 22:11]
  assign io_data_9 = table_9; // @[numa.scala 22:11]
  assign io_data_10 = table_10; // @[numa.scala 22:11]
  assign io_data_11 = table_11; // @[numa.scala 22:11]
  assign io_data_12 = table_12; // @[numa.scala 22:11]
  assign io_data_13 = table_13; // @[numa.scala 22:11]
  assign config_awready = config_wvalid; // @[numa.scala 24:18]
  assign config_arready = ~rvalid; // @[numa.scala 25:28]
  assign config_wready = config_wvalid; // @[numa.scala 23:17]
  assign config_rdata = 5'h1f == eraddr ? table_31 : _GEN_671; // @[numa.scala 76:16 numa.scala 76:16]
  assign config_rvalid = rvalid; // @[numa.scala 26:17]
  assign config_bvalid = bvalid; // @[numa.scala 27:17]
  always @(posedge clock) begin
    if (reset) begin // @[numa.scala 17:22]
      table_0 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h0 == io_wptr_1) begin // @[numa.scala 46:23]
        table_0 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_0 <= _GEN_64;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_0 <= _GEN_64;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_0 <= _GEN_224;
    end else begin
      table_0 <= _GEN_512;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_1 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h1 == io_wptr_1) begin // @[numa.scala 46:23]
        table_1 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_1 <= _GEN_65;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_1 <= _GEN_65;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_1 <= _GEN_225;
    end else begin
      table_1 <= _GEN_513;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_2 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h2 == io_wptr_1) begin // @[numa.scala 46:23]
        table_2 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_2 <= _GEN_66;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_2 <= _GEN_66;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_2 <= _GEN_226;
    end else begin
      table_2 <= _GEN_514;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_3 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h3 == io_wptr_1) begin // @[numa.scala 46:23]
        table_3 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_3 <= _GEN_67;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_3 <= _GEN_67;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_3 <= _GEN_227;
    end else begin
      table_3 <= _GEN_515;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_4 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h4 == io_wptr_1) begin // @[numa.scala 46:23]
        table_4 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_4 <= _GEN_68;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_4 <= _GEN_68;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_4 <= _GEN_228;
    end else begin
      table_4 <= _GEN_516;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_5 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h5 == io_wptr_1) begin // @[numa.scala 46:23]
        table_5 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_5 <= _GEN_69;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_5 <= _GEN_69;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_5 <= _GEN_229;
    end else begin
      table_5 <= _GEN_517;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_6 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h6 == io_wptr_1) begin // @[numa.scala 46:23]
        table_6 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_6 <= _GEN_70;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_6 <= _GEN_70;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_6 <= _GEN_230;
    end else begin
      table_6 <= _GEN_518;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_7 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h7 == io_wptr_1) begin // @[numa.scala 46:23]
        table_7 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_7 <= _GEN_71;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_7 <= _GEN_71;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_7 <= _GEN_231;
    end else begin
      table_7 <= _GEN_519;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_8 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h8 == io_wptr_1) begin // @[numa.scala 46:23]
        table_8 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_8 <= _GEN_72;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_8 <= _GEN_72;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_8 <= _GEN_232;
    end else begin
      table_8 <= _GEN_520;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_9 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h9 == io_wptr_1) begin // @[numa.scala 46:23]
        table_9 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_9 <= _GEN_73;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_9 <= _GEN_73;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_9 <= _GEN_233;
    end else begin
      table_9 <= _GEN_521;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_10 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'ha == io_wptr_1) begin // @[numa.scala 46:23]
        table_10 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_10 <= _GEN_74;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_10 <= _GEN_74;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_10 <= _GEN_234;
    end else begin
      table_10 <= _GEN_522;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_11 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'hb == io_wptr_1) begin // @[numa.scala 46:23]
        table_11 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_11 <= _GEN_75;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_11 <= _GEN_75;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_11 <= _GEN_235;
    end else begin
      table_11 <= _GEN_523;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_12 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'hc == io_wptr_1) begin // @[numa.scala 46:23]
        table_12 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_12 <= _GEN_76;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_12 <= _GEN_76;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_12 <= _GEN_236;
    end else begin
      table_12 <= _GEN_524;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_13 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'hd == io_wptr_1) begin // @[numa.scala 46:23]
        table_13 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_13 <= _GEN_77;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_13 <= _GEN_77;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_13 <= _GEN_237;
    end else begin
      table_13 <= _GEN_525;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_14 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'he == io_wptr_1) begin // @[numa.scala 46:23]
        table_14 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_14 <= _GEN_78;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_14 <= _GEN_78;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_14 <= _GEN_238;
    end else begin
      table_14 <= _GEN_526;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_15 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'hf == io_wptr_1) begin // @[numa.scala 46:23]
        table_15 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_15 <= _GEN_79;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_15 <= _GEN_79;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_15 <= _GEN_239;
    end else begin
      table_15 <= _GEN_527;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_16 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h10 == io_wptr_1) begin // @[numa.scala 46:23]
        table_16 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_16 <= _GEN_80;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_16 <= _GEN_80;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_16 <= _GEN_240;
    end else begin
      table_16 <= _GEN_528;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_17 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h11 == io_wptr_1) begin // @[numa.scala 46:23]
        table_17 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_17 <= _GEN_81;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_17 <= _GEN_81;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_17 <= _GEN_241;
    end else begin
      table_17 <= _GEN_529;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_18 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h12 == io_wptr_1) begin // @[numa.scala 46:23]
        table_18 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_18 <= _GEN_82;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_18 <= _GEN_82;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_18 <= _GEN_242;
    end else begin
      table_18 <= _GEN_530;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_19 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h13 == io_wptr_1) begin // @[numa.scala 46:23]
        table_19 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_19 <= _GEN_83;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_19 <= _GEN_83;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_19 <= _GEN_243;
    end else begin
      table_19 <= _GEN_531;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_20 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h14 == io_wptr_1) begin // @[numa.scala 46:23]
        table_20 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_20 <= _GEN_84;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_20 <= _GEN_84;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_20 <= _GEN_244;
    end else begin
      table_20 <= _GEN_532;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_21 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h15 == io_wptr_1) begin // @[numa.scala 46:23]
        table_21 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_21 <= _GEN_85;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_21 <= _GEN_85;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_21 <= _GEN_245;
    end else begin
      table_21 <= _GEN_533;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_22 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h16 == io_wptr_1) begin // @[numa.scala 46:23]
        table_22 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_22 <= _GEN_86;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_22 <= _GEN_86;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_22 <= _GEN_246;
    end else begin
      table_22 <= _GEN_534;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_23 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h17 == io_wptr_1) begin // @[numa.scala 46:23]
        table_23 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_23 <= _GEN_87;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_23 <= _GEN_87;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_23 <= _GEN_247;
    end else begin
      table_23 <= _GEN_535;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_24 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h18 == io_wptr_1) begin // @[numa.scala 46:23]
        table_24 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_24 <= _GEN_88;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_24 <= _GEN_88;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_24 <= _GEN_248;
    end else begin
      table_24 <= _GEN_536;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_25 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h19 == io_wptr_1) begin // @[numa.scala 46:23]
        table_25 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_25 <= _GEN_89;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_25 <= _GEN_89;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_25 <= _GEN_249;
    end else begin
      table_25 <= _GEN_537;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_26 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h1a == io_wptr_1) begin // @[numa.scala 46:23]
        table_26 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_26 <= _GEN_90;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_26 <= _GEN_90;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_26 <= _GEN_250;
    end else begin
      table_26 <= _GEN_538;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_27 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h1b == io_wptr_1) begin // @[numa.scala 46:23]
        table_27 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_27 <= _GEN_91;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_27 <= _GEN_91;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_27 <= _GEN_251;
    end else begin
      table_27 <= _GEN_539;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_28 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h1c == io_wptr_1) begin // @[numa.scala 46:23]
        table_28 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_28 <= _GEN_92;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_28 <= _GEN_92;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_28 <= _GEN_252;
    end else begin
      table_28 <= _GEN_540;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_29 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h1d == io_wptr_1) begin // @[numa.scala 46:23]
        table_29 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_29 <= _GEN_93;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_29 <= _GEN_93;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_29 <= _GEN_253;
    end else begin
      table_29 <= _GEN_541;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_30 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h1e == io_wptr_1) begin // @[numa.scala 46:23]
        table_30 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_30 <= _GEN_94;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_30 <= _GEN_94;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_30 <= _GEN_254;
    end else begin
      table_30 <= _GEN_542;
    end
    if (reset) begin // @[numa.scala 17:22]
      table_31 <= 32'h0; // @[numa.scala 17:22]
    end else if (config_wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[numa.scala 43:50]
      if (5'h1f == io_wptr_1) begin // @[numa.scala 46:23]
        table_31 <= io_dataIn_1; // @[numa.scala 46:23]
      end else begin
        table_31 <= _GEN_95;
      end
    end else if (config_wvalid & io_writeFlag_0) begin // @[numa.scala 47:47]
      table_31 <= _GEN_95;
    end else if (config_wvalid & io_writeFlag_1) begin // @[numa.scala 50:47]
      table_31 <= _GEN_255;
    end else begin
      table_31 <= _GEN_543;
    end
    if (reset) begin // @[numa.scala 18:23]
      rvalid <= 1'h0; // @[numa.scala 18:23]
    end else begin
      rvalid <= _GEN_674;
    end
    if (reset) begin // @[numa.scala 19:23]
      bvalid <= 1'h0; // @[numa.scala 19:23]
    end else begin
      bvalid <= _GEN_676;
    end
    if (config_arvalid & config_arready) begin // @[numa.scala 69:41]
      eraddr <= config_araddr[6:2]; // @[numa.scala 70:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  table_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  table_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  table_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  table_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  table_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  table_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  table_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  table_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  table_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  table_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  table_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  table_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  table_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  table_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  table_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  table_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  table_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  table_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  table_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  table_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  table_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  table_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  table_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  table_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  table_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  table_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  table_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  table_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  table_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  table_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  table_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  table_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  rvalid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  bvalid = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  eraddr = _RAND_34[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module controller(
  input         clock,
  input         reset,
  output [31:0] io_data_0,
  output [31:0] io_data_1,
  output [31:0] io_data_2,
  output [31:0] io_data_3,
  output [31:0] io_data_4,
  output [31:0] io_data_5,
  output [31:0] io_data_6,
  output [31:0] io_data_7,
  output [31:0] io_data_8,
  output [31:0] io_data_9,
  output [31:0] io_data_10,
  output [31:0] io_data_11,
  input         io_fin_0,
  input         io_fin_1,
  input         io_fin_2,
  input         io_fin_3,
  input         io_fin_4,
  input         io_fin_5,
  input         io_fin_6,
  input         io_fin_7,
  input         io_fin_8,
  input         io_fin_9,
  input         io_fin_10,
  input         io_fin_11,
  input         io_fin_12,
  input         io_fin_13,
  input         io_fin_14,
  input         io_fin_15,
  output        io_signal,
  output        io_start,
  output [31:0] io_level,
  input  [31:0] io_unvisited_size,
  input  [63:0] io_traveled_edges,
  input  [63:0] io_config_awaddr,
  output        io_config_awready,
  input  [63:0] io_config_araddr,
  input         io_config_arvalid,
  output        io_config_arready,
  input  [31:0] io_config_wdata,
  input  [3:0]  io_config_wstrb,
  input         io_config_wvalid,
  output        io_config_wready,
  output [31:0] io_config_rdata,
  output        io_config_rvalid,
  input         io_config_rready,
  output        io_config_bvalid,
  input         io_config_bready,
  output        io_flush_cache,
  input         io_flush_cache_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  controls_clock; // @[BFS.scala 1098:24]
  wire  controls_reset; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_0; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_1; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_2; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_3; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_4; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_5; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_6; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_7; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_8; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_9; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_10; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_11; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_12; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_data_13; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_dataIn_0; // @[BFS.scala 1098:24]
  wire [31:0] controls_io_dataIn_1; // @[BFS.scala 1098:24]
  wire  controls_io_writeFlag_0; // @[BFS.scala 1098:24]
  wire  controls_io_writeFlag_1; // @[BFS.scala 1098:24]
  wire [4:0] controls_io_wptr_0; // @[BFS.scala 1098:24]
  wire [4:0] controls_io_wptr_1; // @[BFS.scala 1098:24]
  wire [63:0] controls_config_awaddr; // @[BFS.scala 1098:24]
  wire  controls_config_awready; // @[BFS.scala 1098:24]
  wire [63:0] controls_config_araddr; // @[BFS.scala 1098:24]
  wire  controls_config_arvalid; // @[BFS.scala 1098:24]
  wire  controls_config_arready; // @[BFS.scala 1098:24]
  wire [31:0] controls_config_wdata; // @[BFS.scala 1098:24]
  wire [3:0] controls_config_wstrb; // @[BFS.scala 1098:24]
  wire  controls_config_wvalid; // @[BFS.scala 1098:24]
  wire  controls_config_wready; // @[BFS.scala 1098:24]
  wire [31:0] controls_config_rdata; // @[BFS.scala 1098:24]
  wire  controls_config_rvalid; // @[BFS.scala 1098:24]
  wire  controls_config_rready; // @[BFS.scala 1098:24]
  wire  controls_config_bvalid; // @[BFS.scala 1098:24]
  wire  controls_config_bready; // @[BFS.scala 1098:24]
  reg [31:0] level; // @[BFS.scala 1099:22]
  reg [2:0] status; // @[BFS.scala 1109:23]
  wire  start = controls_io_data_0[0]; // @[BFS.scala 1110:34]
  reg  FIN_0; // @[BFS.scala 1111:20]
  reg  FIN_1; // @[BFS.scala 1111:20]
  reg  FIN_2; // @[BFS.scala 1111:20]
  reg  FIN_3; // @[BFS.scala 1111:20]
  reg  FIN_4; // @[BFS.scala 1111:20]
  reg  FIN_5; // @[BFS.scala 1111:20]
  reg  FIN_6; // @[BFS.scala 1111:20]
  reg  FIN_7; // @[BFS.scala 1111:20]
  reg  FIN_8; // @[BFS.scala 1111:20]
  reg  FIN_9; // @[BFS.scala 1111:20]
  reg  FIN_10; // @[BFS.scala 1111:20]
  reg  FIN_11; // @[BFS.scala 1111:20]
  reg  FIN_12; // @[BFS.scala 1111:20]
  reg  FIN_13; // @[BFS.scala 1111:20]
  reg  FIN_14; // @[BFS.scala 1111:20]
  reg  FIN_15; // @[BFS.scala 1111:20]
  wire [63:0] _new_tep_T = {controls_io_data_12,controls_io_data_13}; // @[Cat.scala 30:58]
  wire [63:0] new_tep = _new_tep_T + io_traveled_edges; // @[BFS.scala 1112:65]
  reg [63:0] counterValue; // @[BFS.scala 1113:29]
  wire  _controls_io_writeFlag_0_T = status == 3'h3; // @[BFS.scala 1116:38]
  wire  _controls_io_writeFlag_0_T_1 = status == 3'h2; // @[BFS.scala 1116:58]
  wire  _controls_io_writeFlag_0_T_3 = status == 3'h6; // @[BFS.scala 1116:78]
  wire [3:0] _controls_io_wptr_0_T_3 = _controls_io_writeFlag_0_T_1 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_0_T_4 = _controls_io_writeFlag_0_T_3 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_0_T_6 = _controls_io_wptr_0_T_3 | _controls_io_wptr_0_T_4; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_5 = _controls_io_writeFlag_0_T_1 ? new_tep[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_6 = _controls_io_writeFlag_0_T_3 ? counterValue[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [1:0] _controls_io_dataIn_0_T_7 = _controls_io_writeFlag_0_T ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_8 = _controls_io_dataIn_0_T_5 | _controls_io_dataIn_0_T_6; // @[Mux.scala 27:72]
  wire [31:0] _GEN_43 = {{30'd0}, _controls_io_dataIn_0_T_7}; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_1_T_1 = _controls_io_writeFlag_0_T_1 ? 4'hd : 4'hf; // @[BFS.scala 1128:29]
  wire [31:0] _controls_io_dataIn_1_T_4 = _controls_io_writeFlag_0_T_1 ? new_tep[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_1_T_5 = _controls_io_writeFlag_0_T_3 ? counterValue[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1 = status == 3'h0 & start; // @[BFS.scala 1134:28]
  wire  _T_2 = status == 3'h4; // @[BFS.scala 1136:21]
  wire [2:0] _GEN_0 = io_unvisited_size == 32'h0 ? 3'h6 : 3'h1; // @[BFS.scala 1141:36 BFS.scala 1142:14 BFS.scala 1144:14]
  wire [2:0] _GEN_1 = _controls_io_writeFlag_0_T ? 3'h0 : status; // @[BFS.scala 1150:32 BFS.scala 1151:12 BFS.scala 1109:23]
  wire [2:0] _GEN_2 = _controls_io_writeFlag_0_T_3 ? 3'h5 : _GEN_1; // @[BFS.scala 1148:40 BFS.scala 1149:12]
  wire [2:0] _GEN_3 = status == 3'h5 & io_flush_cache_end ? 3'h3 : _GEN_2; // @[BFS.scala 1146:62 BFS.scala 1147:12]
  wire [2:0] _GEN_4 = _controls_io_writeFlag_0_T_1 ? _GEN_0 : _GEN_3; // @[BFS.scala 1140:32]
  wire  _GEN_8 = io_signal ? 1'h0 : FIN_0; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_9 = io_fin_0 | _GEN_8; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_10 = io_signal ? 1'h0 : FIN_1; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_11 = io_fin_1 | _GEN_10; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_12 = io_signal ? 1'h0 : FIN_2; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_13 = io_fin_2 | _GEN_12; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_14 = io_signal ? 1'h0 : FIN_3; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_15 = io_fin_3 | _GEN_14; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_16 = io_signal ? 1'h0 : FIN_4; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_17 = io_fin_4 | _GEN_16; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_18 = io_signal ? 1'h0 : FIN_5; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_19 = io_fin_5 | _GEN_18; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_20 = io_signal ? 1'h0 : FIN_6; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_21 = io_fin_6 | _GEN_20; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_22 = io_signal ? 1'h0 : FIN_7; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_23 = io_fin_7 | _GEN_22; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_24 = io_signal ? 1'h0 : FIN_8; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_25 = io_fin_8 | _GEN_24; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_26 = io_signal ? 1'h0 : FIN_9; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_27 = io_fin_9 | _GEN_26; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_28 = io_signal ? 1'h0 : FIN_10; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_29 = io_fin_10 | _GEN_28; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_30 = io_signal ? 1'h0 : FIN_11; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_31 = io_fin_11 | _GEN_30; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_32 = io_signal ? 1'h0 : FIN_12; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_33 = io_fin_12 | _GEN_32; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_34 = io_signal ? 1'h0 : FIN_13; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_35 = io_fin_13 | _GEN_34; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_36 = io_signal ? 1'h0 : FIN_14; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_37 = io_fin_14 | _GEN_36; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire  _GEN_38 = io_signal ? 1'h0 : FIN_15; // @[BFS.scala 1158:28 BFS.scala 1159:11 BFS.scala 1111:20]
  wire  _GEN_39 = io_fin_15 | _GEN_38; // @[BFS.scala 1156:22 BFS.scala 1157:11]
  wire [31:0] _level_T_1 = level + 32'h1; // @[BFS.scala 1165:20]
  wire [63:0] _counterValue_T_1 = counterValue + 64'h1; // @[BFS.scala 1173:34]
  LookupTable controls ( // @[BFS.scala 1098:24]
    .clock(controls_clock),
    .reset(controls_reset),
    .io_data_0(controls_io_data_0),
    .io_data_1(controls_io_data_1),
    .io_data_2(controls_io_data_2),
    .io_data_3(controls_io_data_3),
    .io_data_4(controls_io_data_4),
    .io_data_5(controls_io_data_5),
    .io_data_6(controls_io_data_6),
    .io_data_7(controls_io_data_7),
    .io_data_8(controls_io_data_8),
    .io_data_9(controls_io_data_9),
    .io_data_10(controls_io_data_10),
    .io_data_11(controls_io_data_11),
    .io_data_12(controls_io_data_12),
    .io_data_13(controls_io_data_13),
    .io_dataIn_0(controls_io_dataIn_0),
    .io_dataIn_1(controls_io_dataIn_1),
    .io_writeFlag_0(controls_io_writeFlag_0),
    .io_writeFlag_1(controls_io_writeFlag_1),
    .io_wptr_0(controls_io_wptr_0),
    .io_wptr_1(controls_io_wptr_1),
    .config_awaddr(controls_config_awaddr),
    .config_awready(controls_config_awready),
    .config_araddr(controls_config_araddr),
    .config_arvalid(controls_config_arvalid),
    .config_arready(controls_config_arready),
    .config_wdata(controls_config_wdata),
    .config_wstrb(controls_config_wstrb),
    .config_wvalid(controls_config_wvalid),
    .config_wready(controls_config_wready),
    .config_rdata(controls_config_rdata),
    .config_rvalid(controls_config_rvalid),
    .config_rready(controls_config_rready),
    .config_bvalid(controls_config_bvalid),
    .config_bready(controls_config_bready)
  );
  assign io_data_0 = controls_io_data_0; // @[BFS.scala 1177:11]
  assign io_data_1 = controls_io_data_1; // @[BFS.scala 1177:11]
  assign io_data_2 = controls_io_data_2; // @[BFS.scala 1177:11]
  assign io_data_3 = controls_io_data_3; // @[BFS.scala 1177:11]
  assign io_data_4 = controls_io_data_4; // @[BFS.scala 1177:11]
  assign io_data_5 = controls_io_data_5; // @[BFS.scala 1177:11]
  assign io_data_6 = controls_io_data_6; // @[BFS.scala 1177:11]
  assign io_data_7 = controls_io_data_7; // @[BFS.scala 1177:11]
  assign io_data_8 = controls_io_data_8; // @[BFS.scala 1177:11]
  assign io_data_9 = controls_io_data_9; // @[BFS.scala 1177:11]
  assign io_data_10 = controls_io_data_10; // @[BFS.scala 1177:11]
  assign io_data_11 = controls_io_data_11; // @[BFS.scala 1177:11]
  assign io_signal = _T_2 | _controls_io_writeFlag_0_T_1; // @[BFS.scala 1176:36]
  assign io_start = status == 3'h4; // @[BFS.scala 1179:22]
  assign io_level = level; // @[BFS.scala 1178:12]
  assign io_config_awready = controls_config_awready; // @[BFS.scala 1115:19]
  assign io_config_arready = controls_config_arready; // @[BFS.scala 1115:19]
  assign io_config_wready = controls_config_wready; // @[BFS.scala 1115:19]
  assign io_config_rdata = controls_config_rdata; // @[BFS.scala 1115:19]
  assign io_config_rvalid = controls_config_rvalid; // @[BFS.scala 1115:19]
  assign io_config_bvalid = controls_config_bvalid; // @[BFS.scala 1115:19]
  assign io_flush_cache = status == 3'h5; // @[BFS.scala 1180:28]
  assign controls_clock = clock;
  assign controls_reset = reset;
  assign controls_io_dataIn_0 = _controls_io_dataIn_0_T_8 | _GEN_43; // @[Mux.scala 27:72]
  assign controls_io_dataIn_1 = _controls_io_dataIn_1_T_4 | _controls_io_dataIn_1_T_5; // @[Mux.scala 27:72]
  assign controls_io_writeFlag_0 = status == 3'h3 | status == 3'h2 | status == 3'h6; // @[BFS.scala 1116:69]
  assign controls_io_writeFlag_1 = _controls_io_writeFlag_0_T_1 | _controls_io_writeFlag_0_T_3; // @[BFS.scala 1127:49]
  assign controls_io_wptr_0 = {{1'd0}, _controls_io_wptr_0_T_6}; // @[Mux.scala 27:72]
  assign controls_io_wptr_1 = {{1'd0}, _controls_io_wptr_1_T_1}; // @[BFS.scala 1128:29]
  assign controls_config_awaddr = io_config_awaddr; // @[BFS.scala 1115:19]
  assign controls_config_araddr = io_config_araddr; // @[BFS.scala 1115:19]
  assign controls_config_arvalid = io_config_arvalid; // @[BFS.scala 1115:19]
  assign controls_config_wdata = io_config_wdata; // @[BFS.scala 1115:19]
  assign controls_config_wstrb = io_config_wstrb; // @[BFS.scala 1115:19]
  assign controls_config_wvalid = io_config_wvalid; // @[BFS.scala 1115:19]
  assign controls_config_rready = io_config_rready; // @[BFS.scala 1115:19]
  assign controls_config_bready = io_config_bready; // @[BFS.scala 1115:19]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1099:22]
      level <= 32'h0; // @[BFS.scala 1099:22]
    end else if (_controls_io_writeFlag_0_T_1) begin // @[BFS.scala 1164:26]
      level <= _level_T_1; // @[BFS.scala 1165:11]
    end else if (_T_1) begin // @[BFS.scala 1166:43]
      level <= 32'hffffffff; // @[BFS.scala 1167:11]
    end
    if (reset) begin // @[BFS.scala 1109:23]
      status <= 3'h0; // @[BFS.scala 1109:23]
    end else if (status == 3'h0 & start) begin // @[BFS.scala 1134:37]
      status <= 3'h4; // @[BFS.scala 1135:12]
    end else if (status == 3'h4) begin // @[BFS.scala 1136:34]
      status <= 3'h1; // @[BFS.scala 1137:12]
    end else if (status == 3'h1 & (FIN_0 & FIN_1 & FIN_2 & FIN_3 & FIN_4 & FIN_5 & FIN_6 & FIN_7 & FIN_8 & FIN_9 &
      FIN_10 & FIN_11 & FIN_12 & FIN_13 & FIN_14 & FIN_15)) begin // @[BFS.scala 1138:51]
      status <= 3'h2; // @[BFS.scala 1139:12]
    end else begin
      status <= _GEN_4;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_0 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_0 <= _GEN_9;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_1 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_1 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_2 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_2 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_3 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_3 <= _GEN_15;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_4 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_4 <= _GEN_17;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_5 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_5 <= _GEN_19;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_6 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_6 <= _GEN_21;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_7 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_7 <= _GEN_23;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_8 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_8 <= _GEN_25;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_9 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_9 <= _GEN_27;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_10 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_10 <= _GEN_29;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_11 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_11 <= _GEN_31;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_12 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_12 <= _GEN_33;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_13 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_13 <= _GEN_35;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_14 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_14 <= _GEN_37;
    end
    if (reset) begin // @[BFS.scala 1111:20]
      FIN_15 <= 1'h0; // @[BFS.scala 1111:20]
    end else begin
      FIN_15 <= _GEN_39;
    end
    if (reset) begin // @[BFS.scala 1113:29]
      counterValue <= 64'h0; // @[BFS.scala 1113:29]
    end else if (_T_2) begin // @[BFS.scala 1170:29]
      counterValue <= 64'h0; // @[BFS.scala 1171:18]
    end else begin
      counterValue <= _counterValue_T_1; // @[BFS.scala 1173:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  level = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  status = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  FIN_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIN_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  FIN_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  FIN_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  FIN_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  FIN_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  FIN_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  FIN_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  FIN_8 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  FIN_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  FIN_10 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  FIN_11 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  FIN_12 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  FIN_13 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  FIN_14 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  FIN_15 = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  counterValue = _RAND_18[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pipeline(
  input         clock,
  input         reset,
  input         io_dout_ready,
  output        io_dout_valid,
  output [31:0] io_dout_bits_tdata,
  output        io_din_ready,
  input         io_din_valid,
  input  [31:0] io_din_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] data_tdata; // @[util.scala 143:21]
  reg  valid; // @[util.scala 144:22]
  assign io_dout_valid = valid; // @[util.scala 151:17]
  assign io_dout_bits_tdata = data_tdata; // @[util.scala 152:16]
  assign io_din_ready = io_dout_ready; // @[util.scala 150:16]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 143:21]
      data_tdata <= 32'h0; // @[util.scala 143:21]
    end else if (io_dout_ready) begin // @[util.scala 145:22]
      data_tdata <= io_din_bits_tdata; // @[util.scala 146:10]
    end
    if (reset) begin // @[util.scala 144:22]
      valid <= 1'h0; // @[util.scala 144:22]
    end else if (io_dout_ready) begin // @[util.scala 145:22]
      valid <= io_din_valid; // @[util.scala 147:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_tdata = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  valid = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multi_channel_fifo(
  input          clock,
  input          reset,
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [31:0]  io_in_0_bits_tdata,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [31:0]  io_in_1_bits_tdata,
  output         io_in_2_ready,
  input          io_in_2_valid,
  input  [31:0]  io_in_2_bits_tdata,
  output         io_in_3_ready,
  input          io_in_3_valid,
  input  [31:0]  io_in_3_bits_tdata,
  output         io_in_4_ready,
  input          io_in_4_valid,
  input  [31:0]  io_in_4_bits_tdata,
  output         io_in_5_ready,
  input          io_in_5_valid,
  input  [31:0]  io_in_5_bits_tdata,
  output         io_in_6_ready,
  input          io_in_6_valid,
  input  [31:0]  io_in_6_bits_tdata,
  output         io_in_7_ready,
  input          io_in_7_valid,
  input  [31:0]  io_in_7_bits_tdata,
  output         io_in_8_ready,
  input          io_in_8_valid,
  input  [31:0]  io_in_8_bits_tdata,
  output         io_in_9_ready,
  input          io_in_9_valid,
  input  [31:0]  io_in_9_bits_tdata,
  output         io_in_10_ready,
  input          io_in_10_valid,
  input  [31:0]  io_in_10_bits_tdata,
  output         io_in_11_ready,
  input          io_in_11_valid,
  input  [31:0]  io_in_11_bits_tdata,
  output         io_in_12_ready,
  input          io_in_12_valid,
  input  [31:0]  io_in_12_bits_tdata,
  output         io_in_13_ready,
  input          io_in_13_valid,
  input  [31:0]  io_in_13_bits_tdata,
  output         io_in_14_ready,
  input          io_in_14_valid,
  input  [31:0]  io_in_14_bits_tdata,
  output         io_in_15_ready,
  input          io_in_15_valid,
  input  [31:0]  io_in_15_bits_tdata,
  output         io_out_full,
  input  [511:0] io_out_din,
  input          io_out_wr_en,
  output [511:0] io_out_dout,
  input          io_out_rd_en,
  output [8:0]   io_out_data_count,
  output         io_out_valid,
  input          io_flush,
  input          io_is_current_tier
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  collector_fifos_0_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_0_din; // @[BFS.scala 826:16]
  wire  collector_fifos_0_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_0_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_0_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_0_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_0_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_0_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_0_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_0_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_1_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_1_din; // @[BFS.scala 826:16]
  wire  collector_fifos_1_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_1_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_1_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_1_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_1_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_1_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_1_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_1_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_2_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_2_din; // @[BFS.scala 826:16]
  wire  collector_fifos_2_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_2_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_2_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_2_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_2_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_2_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_2_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_2_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_3_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_3_din; // @[BFS.scala 826:16]
  wire  collector_fifos_3_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_3_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_3_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_3_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_3_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_3_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_3_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_3_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_4_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_4_din; // @[BFS.scala 826:16]
  wire  collector_fifos_4_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_4_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_4_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_4_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_4_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_4_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_4_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_4_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_5_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_5_din; // @[BFS.scala 826:16]
  wire  collector_fifos_5_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_5_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_5_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_5_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_5_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_5_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_5_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_5_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_6_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_6_din; // @[BFS.scala 826:16]
  wire  collector_fifos_6_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_6_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_6_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_6_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_6_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_6_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_6_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_6_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_7_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_7_din; // @[BFS.scala 826:16]
  wire  collector_fifos_7_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_7_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_7_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_7_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_7_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_7_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_7_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_7_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_8_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_8_din; // @[BFS.scala 826:16]
  wire  collector_fifos_8_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_8_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_8_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_8_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_8_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_8_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_8_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_8_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_9_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_9_din; // @[BFS.scala 826:16]
  wire  collector_fifos_9_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_9_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_9_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_9_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_9_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_9_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_9_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_9_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_10_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_10_din; // @[BFS.scala 826:16]
  wire  collector_fifos_10_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_10_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_10_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_10_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_10_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_10_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_10_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_10_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_11_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_11_din; // @[BFS.scala 826:16]
  wire  collector_fifos_11_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_11_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_11_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_11_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_11_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_11_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_11_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_11_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_12_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_12_din; // @[BFS.scala 826:16]
  wire  collector_fifos_12_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_12_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_12_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_12_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_12_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_12_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_12_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_12_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_13_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_13_din; // @[BFS.scala 826:16]
  wire  collector_fifos_13_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_13_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_13_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_13_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_13_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_13_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_13_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_13_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_14_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_14_din; // @[BFS.scala 826:16]
  wire  collector_fifos_14_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_14_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_14_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_14_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_14_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_14_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_14_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_14_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_15_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_15_din; // @[BFS.scala 826:16]
  wire  collector_fifos_15_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_15_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_15_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_15_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_15_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_15_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_15_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_15_valid; // @[BFS.scala 826:16]
  wire  in_pipeline_0_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_0_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_0_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_0_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_0_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_0_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_0_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_0_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_1_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_1_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_1_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_1_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_1_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_1_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_1_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_1_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_2_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_2_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_2_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_2_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_2_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_2_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_2_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_2_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_3_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_3_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_3_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_3_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_3_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_3_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_3_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_3_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_4_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_4_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_4_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_4_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_4_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_4_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_4_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_4_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_5_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_5_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_5_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_5_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_5_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_5_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_5_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_5_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_6_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_6_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_6_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_6_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_6_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_6_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_6_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_6_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_7_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_7_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_7_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_7_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_7_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_7_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_7_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_7_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_8_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_8_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_8_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_8_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_8_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_8_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_8_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_8_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_9_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_9_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_9_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_9_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_9_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_9_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_9_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_9_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_10_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_10_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_10_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_10_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_10_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_10_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_10_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_10_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_11_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_11_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_11_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_11_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_11_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_11_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_11_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_11_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_12_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_12_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_12_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_12_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_12_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_12_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_12_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_12_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_13_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_13_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_13_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_13_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_13_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_13_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_13_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_13_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_14_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_14_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_14_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_14_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_14_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_14_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_14_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_14_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_15_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_15_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_15_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_15_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_15_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_15_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_15_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_15_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  _fifos_ready_T_15 = ~collector_fifos_15_full; // @[BFS.scala 828:70]
  wire  fifos_ready = ~collector_fifos_0_full & ~collector_fifos_1_full & ~collector_fifos_2_full & ~
    collector_fifos_3_full & ~collector_fifos_4_full & ~collector_fifos_5_full & ~collector_fifos_6_full & ~
    collector_fifos_7_full & ~collector_fifos_8_full & ~collector_fifos_9_full & ~collector_fifos_10_full & ~
    collector_fifos_11_full & ~collector_fifos_12_full & ~collector_fifos_13_full & ~collector_fifos_14_full &
    _fifos_ready_T_15; // @[BFS.scala 828:91]
  reg [3:0] counter; // @[BFS.scala 829:24]
  wire  _steps_T = in_pipeline_0_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire  _steps_T_2 = in_pipeline_1_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE = {{4'd0}, _steps_T}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] _steps_WIRE_1 = {{4'd0}, _steps_T_2}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_1 = _steps_WIRE + _steps_WIRE_1; // @[BFS.scala 842:107]
  wire  _steps_T_6 = in_pipeline_2_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_4 = {{4'd0}, _steps_T_6}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_2 = steps_1 + _steps_WIRE_4; // @[BFS.scala 842:107]
  wire  _steps_T_13 = in_pipeline_3_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_8 = {{4'd0}, _steps_T_13}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_3 = steps_2 + _steps_WIRE_8; // @[BFS.scala 842:107]
  wire  _steps_T_23 = in_pipeline_4_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_13 = {{4'd0}, _steps_T_23}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_4 = steps_3 + _steps_WIRE_13; // @[BFS.scala 842:107]
  wire  _steps_T_36 = in_pipeline_5_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_19 = {{4'd0}, _steps_T_36}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_5 = steps_4 + _steps_WIRE_19; // @[BFS.scala 842:107]
  wire  _steps_T_52 = in_pipeline_6_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_26 = {{4'd0}, _steps_T_52}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_6 = steps_5 + _steps_WIRE_26; // @[BFS.scala 842:107]
  wire  _steps_T_71 = in_pipeline_7_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_34 = {{4'd0}, _steps_T_71}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_7 = steps_6 + _steps_WIRE_34; // @[BFS.scala 842:107]
  wire  _steps_T_93 = in_pipeline_8_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_43 = {{4'd0}, _steps_T_93}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_8 = steps_7 + _steps_WIRE_43; // @[BFS.scala 842:107]
  wire  _steps_T_118 = in_pipeline_9_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_53 = {{4'd0}, _steps_T_118}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_9 = steps_8 + _steps_WIRE_53; // @[BFS.scala 842:107]
  wire  _steps_T_146 = in_pipeline_10_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_64 = {{4'd0}, _steps_T_146}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_10 = steps_9 + _steps_WIRE_64; // @[BFS.scala 842:107]
  wire  _steps_T_177 = in_pipeline_11_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_76 = {{4'd0}, _steps_T_177}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_11 = steps_10 + _steps_WIRE_76; // @[BFS.scala 842:107]
  wire  _steps_T_211 = in_pipeline_12_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_89 = {{4'd0}, _steps_T_211}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_12 = steps_11 + _steps_WIRE_89; // @[BFS.scala 842:107]
  wire  _steps_T_248 = in_pipeline_13_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_103 = {{4'd0}, _steps_T_248}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_13 = steps_12 + _steps_WIRE_103; // @[BFS.scala 842:107]
  wire  _steps_T_288 = in_pipeline_14_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_118 = {{4'd0}, _steps_T_288}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_14 = steps_13 + _steps_WIRE_118; // @[BFS.scala 842:107]
  wire  _steps_T_331 = in_pipeline_15_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_134 = {{4'd0}, _steps_T_331}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_15 = steps_14 + _steps_WIRE_134; // @[BFS.scala 842:107]
  wire [4:0] _GEN_2 = {{1'd0}, counter}; // @[BFS.scala 847:15]
  wire [4:0] _counter_T_1 = _GEN_2 + steps_15; // @[BFS.scala 847:15]
  wire [4:0] _counter_T_6 = _counter_T_1 - 5'h10; // @[BFS.scala 847:44]
  wire [4:0] _counter_T_9 = _counter_T_1 >= 5'h10 ? _counter_T_6 : _counter_T_1; // @[BFS.scala 847:8]
  wire [3:0] _GEN_0 = io_flush ? 4'h0 : counter; // @[BFS.scala 855:23 BFS.scala 856:13 BFS.scala 829:24]
  wire [4:0] _GEN_1 = steps_15 != 5'h0 ? _counter_T_9 : {{1'd0}, _GEN_0}; // @[BFS.scala 853:39 BFS.scala 854:13]
  wire [3:0] _fifo_in_data_T_2 = 4'h0 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_4 = 5'h10 - _GEN_2; // @[BFS.scala 850:49]
  wire [5:0] _fifo_in_data_T_5 = {{1'd0}, _fifo_in_data_T_4}; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_7 = counter <= 4'h0 ? {{1'd0}, _fifo_in_data_T_2} : _fifo_in_data_T_5[4:0]; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_9 = _fifo_in_data_T_7 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_10 = _fifo_in_data_T_9 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_21 = _fifo_in_data_T_9 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_32 = _fifo_in_data_T_9 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_43 = _fifo_in_data_T_9 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_54 = _fifo_in_data_T_9 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_65 = _fifo_in_data_T_9 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_76 = _fifo_in_data_T_9 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_87 = _fifo_in_data_T_9 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_98 = _fifo_in_data_T_9 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_109 = _fifo_in_data_T_9 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_120 = _fifo_in_data_T_9 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_131 = _fifo_in_data_T_9 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_142 = _fifo_in_data_T_9 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_153 = _fifo_in_data_T_9 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_164 = _fifo_in_data_T_9 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_175 = _fifo_in_data_T_9 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_176 = _fifo_in_data_T_175 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_177 = _fifo_in_data_T_164 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_176; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_178 = _fifo_in_data_T_153 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_177; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_179 = _fifo_in_data_T_142 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_178; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_180 = _fifo_in_data_T_131 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_179; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_181 = _fifo_in_data_T_120 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_180; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_182 = _fifo_in_data_T_109 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_181; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_183 = _fifo_in_data_T_98 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_182; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_184 = _fifo_in_data_T_87 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_183; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_185 = _fifo_in_data_T_76 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_184; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_186 = _fifo_in_data_T_65 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_185; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_187 = _fifo_in_data_T_54 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_186; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_188 = _fifo_in_data_T_43 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_187; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_189 = _fifo_in_data_T_32 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_188; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_190 = _fifo_in_data_T_21 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_189; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data = _fifo_in_data_T_10 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_190; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_177 = _fifo_in_data_T_164 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_175 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_178 = _fifo_in_data_T_153 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_177; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_179 = _fifo_in_data_T_142 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_178; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_180 = _fifo_in_data_T_131 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_179; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_181 = _fifo_in_data_T_120 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_180; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_182 = _fifo_in_data_T_109 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_181; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_183 = _fifo_in_data_T_98 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_182; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_184 = _fifo_in_data_T_87 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_183; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_185 = _fifo_in_data_T_76 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_184; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_186 = _fifo_in_data_T_65 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_185; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_187 = _fifo_in_data_T_54 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_186; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_188 = _fifo_in_data_T_43 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_187; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_189 = _fifo_in_data_T_32 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_188; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_190 = _fifo_in_data_T_21 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_189; // @[Mux.scala 98:16]
  wire  fifo_in_valid = _fifo_in_data_T_10 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_190; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_193 = 4'h1 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_197 = _fifo_in_data_T_4 + 5'h1; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_198 = counter <= 4'h1 ? {{1'd0}, _fifo_in_data_T_193} : _fifo_in_data_T_197; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_200 = _fifo_in_data_T_198 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_201 = _fifo_in_data_T_200 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_212 = _fifo_in_data_T_200 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_223 = _fifo_in_data_T_200 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_234 = _fifo_in_data_T_200 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_245 = _fifo_in_data_T_200 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_256 = _fifo_in_data_T_200 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_267 = _fifo_in_data_T_200 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_278 = _fifo_in_data_T_200 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_289 = _fifo_in_data_T_200 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_300 = _fifo_in_data_T_200 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_311 = _fifo_in_data_T_200 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_322 = _fifo_in_data_T_200 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_333 = _fifo_in_data_T_200 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_344 = _fifo_in_data_T_200 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_355 = _fifo_in_data_T_200 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_366 = _fifo_in_data_T_200 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_367 = _fifo_in_data_T_366 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_368 = _fifo_in_data_T_355 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_367; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_369 = _fifo_in_data_T_344 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_368; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_370 = _fifo_in_data_T_333 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_369; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_371 = _fifo_in_data_T_322 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_370; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_372 = _fifo_in_data_T_311 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_371; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_373 = _fifo_in_data_T_300 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_372; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_374 = _fifo_in_data_T_289 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_373; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_375 = _fifo_in_data_T_278 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_374; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_376 = _fifo_in_data_T_267 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_375; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_377 = _fifo_in_data_T_256 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_376; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_378 = _fifo_in_data_T_245 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_377; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_379 = _fifo_in_data_T_234 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_378; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_380 = _fifo_in_data_T_223 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_379; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_381 = _fifo_in_data_T_212 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_380; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_1 = _fifo_in_data_T_201 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_381; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_368 = _fifo_in_data_T_355 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_366 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_369 = _fifo_in_data_T_344 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_368; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_370 = _fifo_in_data_T_333 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_369; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_371 = _fifo_in_data_T_322 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_370; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_372 = _fifo_in_data_T_311 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_371; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_373 = _fifo_in_data_T_300 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_372; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_374 = _fifo_in_data_T_289 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_373; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_375 = _fifo_in_data_T_278 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_374; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_376 = _fifo_in_data_T_267 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_375; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_377 = _fifo_in_data_T_256 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_376; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_378 = _fifo_in_data_T_245 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_377; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_379 = _fifo_in_data_T_234 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_378; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_380 = _fifo_in_data_T_223 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_379; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_381 = _fifo_in_data_T_212 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_380; // @[Mux.scala 98:16]
  wire  fifo_in_valid_1 = _fifo_in_data_T_201 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_381; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_384 = 4'h2 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_388 = _fifo_in_data_T_4 + 5'h2; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_389 = counter <= 4'h2 ? {{1'd0}, _fifo_in_data_T_384} : _fifo_in_data_T_388; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_391 = _fifo_in_data_T_389 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_392 = _fifo_in_data_T_391 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_403 = _fifo_in_data_T_391 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_414 = _fifo_in_data_T_391 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_425 = _fifo_in_data_T_391 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_436 = _fifo_in_data_T_391 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_447 = _fifo_in_data_T_391 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_458 = _fifo_in_data_T_391 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_469 = _fifo_in_data_T_391 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_480 = _fifo_in_data_T_391 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_491 = _fifo_in_data_T_391 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_502 = _fifo_in_data_T_391 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_513 = _fifo_in_data_T_391 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_524 = _fifo_in_data_T_391 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_535 = _fifo_in_data_T_391 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_546 = _fifo_in_data_T_391 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_557 = _fifo_in_data_T_391 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_558 = _fifo_in_data_T_557 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_559 = _fifo_in_data_T_546 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_558; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_560 = _fifo_in_data_T_535 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_559; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_561 = _fifo_in_data_T_524 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_560; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_562 = _fifo_in_data_T_513 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_561; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_563 = _fifo_in_data_T_502 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_562; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_564 = _fifo_in_data_T_491 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_563; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_565 = _fifo_in_data_T_480 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_564; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_566 = _fifo_in_data_T_469 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_565; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_567 = _fifo_in_data_T_458 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_566; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_568 = _fifo_in_data_T_447 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_567; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_569 = _fifo_in_data_T_436 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_568; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_570 = _fifo_in_data_T_425 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_569; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_571 = _fifo_in_data_T_414 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_570; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_572 = _fifo_in_data_T_403 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_571; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_2 = _fifo_in_data_T_392 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_572; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_559 = _fifo_in_data_T_546 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_557 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_560 = _fifo_in_data_T_535 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_559; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_561 = _fifo_in_data_T_524 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_560; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_562 = _fifo_in_data_T_513 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_561; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_563 = _fifo_in_data_T_502 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_562; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_564 = _fifo_in_data_T_491 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_563; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_565 = _fifo_in_data_T_480 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_564; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_566 = _fifo_in_data_T_469 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_565; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_567 = _fifo_in_data_T_458 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_566; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_568 = _fifo_in_data_T_447 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_567; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_569 = _fifo_in_data_T_436 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_568; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_570 = _fifo_in_data_T_425 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_569; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_571 = _fifo_in_data_T_414 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_570; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_572 = _fifo_in_data_T_403 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_571; // @[Mux.scala 98:16]
  wire  fifo_in_valid_2 = _fifo_in_data_T_392 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_572; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_575 = 4'h3 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_579 = _fifo_in_data_T_4 + 5'h3; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_580 = counter <= 4'h3 ? {{1'd0}, _fifo_in_data_T_575} : _fifo_in_data_T_579; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_582 = _fifo_in_data_T_580 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_583 = _fifo_in_data_T_582 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_594 = _fifo_in_data_T_582 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_605 = _fifo_in_data_T_582 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_616 = _fifo_in_data_T_582 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_627 = _fifo_in_data_T_582 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_638 = _fifo_in_data_T_582 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_649 = _fifo_in_data_T_582 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_660 = _fifo_in_data_T_582 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_671 = _fifo_in_data_T_582 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_682 = _fifo_in_data_T_582 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_693 = _fifo_in_data_T_582 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_704 = _fifo_in_data_T_582 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_715 = _fifo_in_data_T_582 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_726 = _fifo_in_data_T_582 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_737 = _fifo_in_data_T_582 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_748 = _fifo_in_data_T_582 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_749 = _fifo_in_data_T_748 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_750 = _fifo_in_data_T_737 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_749; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_751 = _fifo_in_data_T_726 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_750; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_752 = _fifo_in_data_T_715 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_751; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_753 = _fifo_in_data_T_704 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_752; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_754 = _fifo_in_data_T_693 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_753; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_755 = _fifo_in_data_T_682 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_754; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_756 = _fifo_in_data_T_671 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_755; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_757 = _fifo_in_data_T_660 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_756; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_758 = _fifo_in_data_T_649 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_757; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_759 = _fifo_in_data_T_638 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_758; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_760 = _fifo_in_data_T_627 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_759; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_761 = _fifo_in_data_T_616 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_760; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_762 = _fifo_in_data_T_605 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_761; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_763 = _fifo_in_data_T_594 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_762; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_3 = _fifo_in_data_T_583 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_763; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_750 = _fifo_in_data_T_737 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_748 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_751 = _fifo_in_data_T_726 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_750; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_752 = _fifo_in_data_T_715 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_751; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_753 = _fifo_in_data_T_704 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_752; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_754 = _fifo_in_data_T_693 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_753; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_755 = _fifo_in_data_T_682 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_754; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_756 = _fifo_in_data_T_671 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_755; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_757 = _fifo_in_data_T_660 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_756; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_758 = _fifo_in_data_T_649 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_757; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_759 = _fifo_in_data_T_638 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_758; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_760 = _fifo_in_data_T_627 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_759; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_761 = _fifo_in_data_T_616 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_760; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_762 = _fifo_in_data_T_605 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_761; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_763 = _fifo_in_data_T_594 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_762; // @[Mux.scala 98:16]
  wire  fifo_in_valid_3 = _fifo_in_data_T_583 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_763; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_766 = 4'h4 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_770 = _fifo_in_data_T_4 + 5'h4; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_771 = counter <= 4'h4 ? {{1'd0}, _fifo_in_data_T_766} : _fifo_in_data_T_770; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_773 = _fifo_in_data_T_771 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_774 = _fifo_in_data_T_773 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_785 = _fifo_in_data_T_773 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_796 = _fifo_in_data_T_773 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_807 = _fifo_in_data_T_773 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_818 = _fifo_in_data_T_773 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_829 = _fifo_in_data_T_773 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_840 = _fifo_in_data_T_773 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_851 = _fifo_in_data_T_773 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_862 = _fifo_in_data_T_773 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_873 = _fifo_in_data_T_773 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_884 = _fifo_in_data_T_773 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_895 = _fifo_in_data_T_773 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_906 = _fifo_in_data_T_773 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_917 = _fifo_in_data_T_773 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_928 = _fifo_in_data_T_773 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_939 = _fifo_in_data_T_773 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_940 = _fifo_in_data_T_939 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_941 = _fifo_in_data_T_928 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_940; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_942 = _fifo_in_data_T_917 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_941; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_943 = _fifo_in_data_T_906 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_942; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_944 = _fifo_in_data_T_895 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_943; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_945 = _fifo_in_data_T_884 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_944; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_946 = _fifo_in_data_T_873 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_945; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_947 = _fifo_in_data_T_862 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_946; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_948 = _fifo_in_data_T_851 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_947; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_949 = _fifo_in_data_T_840 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_948; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_950 = _fifo_in_data_T_829 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_949; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_951 = _fifo_in_data_T_818 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_950; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_952 = _fifo_in_data_T_807 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_951; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_953 = _fifo_in_data_T_796 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_952; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_954 = _fifo_in_data_T_785 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_953; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_4 = _fifo_in_data_T_774 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_954; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_941 = _fifo_in_data_T_928 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_939 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_942 = _fifo_in_data_T_917 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_941; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_943 = _fifo_in_data_T_906 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_942; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_944 = _fifo_in_data_T_895 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_943; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_945 = _fifo_in_data_T_884 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_944; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_946 = _fifo_in_data_T_873 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_945; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_947 = _fifo_in_data_T_862 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_946; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_948 = _fifo_in_data_T_851 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_947; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_949 = _fifo_in_data_T_840 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_948; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_950 = _fifo_in_data_T_829 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_949; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_951 = _fifo_in_data_T_818 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_950; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_952 = _fifo_in_data_T_807 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_951; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_953 = _fifo_in_data_T_796 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_952; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_954 = _fifo_in_data_T_785 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_953; // @[Mux.scala 98:16]
  wire  fifo_in_valid_4 = _fifo_in_data_T_774 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_954; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_957 = 4'h5 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_961 = _fifo_in_data_T_4 + 5'h5; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_962 = counter <= 4'h5 ? {{1'd0}, _fifo_in_data_T_957} : _fifo_in_data_T_961; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_964 = _fifo_in_data_T_962 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_965 = _fifo_in_data_T_964 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_976 = _fifo_in_data_T_964 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_987 = _fifo_in_data_T_964 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_998 = _fifo_in_data_T_964 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1009 = _fifo_in_data_T_964 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1020 = _fifo_in_data_T_964 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1031 = _fifo_in_data_T_964 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1042 = _fifo_in_data_T_964 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1053 = _fifo_in_data_T_964 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1064 = _fifo_in_data_T_964 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1075 = _fifo_in_data_T_964 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1086 = _fifo_in_data_T_964 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1097 = _fifo_in_data_T_964 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1108 = _fifo_in_data_T_964 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1119 = _fifo_in_data_T_964 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1130 = _fifo_in_data_T_964 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1131 = _fifo_in_data_T_1130 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1132 = _fifo_in_data_T_1119 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1131; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1133 = _fifo_in_data_T_1108 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1132; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1134 = _fifo_in_data_T_1097 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1133; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1135 = _fifo_in_data_T_1086 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1134; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1136 = _fifo_in_data_T_1075 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1135; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1137 = _fifo_in_data_T_1064 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1136; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1138 = _fifo_in_data_T_1053 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1137; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1139 = _fifo_in_data_T_1042 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1138; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1140 = _fifo_in_data_T_1031 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1139; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1141 = _fifo_in_data_T_1020 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1140; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1142 = _fifo_in_data_T_1009 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1141; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1143 = _fifo_in_data_T_998 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1142; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1144 = _fifo_in_data_T_987 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1143; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1145 = _fifo_in_data_T_976 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1144; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_5 = _fifo_in_data_T_965 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1145; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1132 = _fifo_in_data_T_1119 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1130 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1133 = _fifo_in_data_T_1108 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1132; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1134 = _fifo_in_data_T_1097 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1133; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1135 = _fifo_in_data_T_1086 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1134; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1136 = _fifo_in_data_T_1075 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1135; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1137 = _fifo_in_data_T_1064 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1136; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1138 = _fifo_in_data_T_1053 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1137; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1139 = _fifo_in_data_T_1042 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1138; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1140 = _fifo_in_data_T_1031 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1139; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1141 = _fifo_in_data_T_1020 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1140; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1142 = _fifo_in_data_T_1009 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1141; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1143 = _fifo_in_data_T_998 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1142; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1144 = _fifo_in_data_T_987 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1143; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1145 = _fifo_in_data_T_976 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1144; // @[Mux.scala 98:16]
  wire  fifo_in_valid_5 = _fifo_in_data_T_965 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1145; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1148 = 4'h6 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1152 = _fifo_in_data_T_4 + 5'h6; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1153 = counter <= 4'h6 ? {{1'd0}, _fifo_in_data_T_1148} : _fifo_in_data_T_1152; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1155 = _fifo_in_data_T_1153 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1156 = _fifo_in_data_T_1155 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1167 = _fifo_in_data_T_1155 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1178 = _fifo_in_data_T_1155 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1189 = _fifo_in_data_T_1155 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1200 = _fifo_in_data_T_1155 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1211 = _fifo_in_data_T_1155 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1222 = _fifo_in_data_T_1155 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1233 = _fifo_in_data_T_1155 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1244 = _fifo_in_data_T_1155 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1255 = _fifo_in_data_T_1155 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1266 = _fifo_in_data_T_1155 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1277 = _fifo_in_data_T_1155 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1288 = _fifo_in_data_T_1155 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1299 = _fifo_in_data_T_1155 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1310 = _fifo_in_data_T_1155 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1321 = _fifo_in_data_T_1155 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1322 = _fifo_in_data_T_1321 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1323 = _fifo_in_data_T_1310 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1322; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1324 = _fifo_in_data_T_1299 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1323; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1325 = _fifo_in_data_T_1288 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1324; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1326 = _fifo_in_data_T_1277 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1325; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1327 = _fifo_in_data_T_1266 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1326; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1328 = _fifo_in_data_T_1255 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1327; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1329 = _fifo_in_data_T_1244 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1328; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1330 = _fifo_in_data_T_1233 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1329; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1331 = _fifo_in_data_T_1222 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1330; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1332 = _fifo_in_data_T_1211 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1331; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1333 = _fifo_in_data_T_1200 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1332; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1334 = _fifo_in_data_T_1189 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1333; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1335 = _fifo_in_data_T_1178 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1334; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1336 = _fifo_in_data_T_1167 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1335; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_6 = _fifo_in_data_T_1156 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1336; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1323 = _fifo_in_data_T_1310 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1321 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1324 = _fifo_in_data_T_1299 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1323; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1325 = _fifo_in_data_T_1288 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1324; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1326 = _fifo_in_data_T_1277 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1325; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1327 = _fifo_in_data_T_1266 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1326; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1328 = _fifo_in_data_T_1255 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1327; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1329 = _fifo_in_data_T_1244 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1328; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1330 = _fifo_in_data_T_1233 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1329; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1331 = _fifo_in_data_T_1222 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1330; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1332 = _fifo_in_data_T_1211 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1331; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1333 = _fifo_in_data_T_1200 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1332; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1334 = _fifo_in_data_T_1189 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1333; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1335 = _fifo_in_data_T_1178 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1334; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1336 = _fifo_in_data_T_1167 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1335; // @[Mux.scala 98:16]
  wire  fifo_in_valid_6 = _fifo_in_data_T_1156 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1336; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1339 = 4'h7 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1343 = _fifo_in_data_T_4 + 5'h7; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1344 = counter <= 4'h7 ? {{1'd0}, _fifo_in_data_T_1339} : _fifo_in_data_T_1343; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1346 = _fifo_in_data_T_1344 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1347 = _fifo_in_data_T_1346 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1358 = _fifo_in_data_T_1346 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1369 = _fifo_in_data_T_1346 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1380 = _fifo_in_data_T_1346 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1391 = _fifo_in_data_T_1346 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1402 = _fifo_in_data_T_1346 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1413 = _fifo_in_data_T_1346 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1424 = _fifo_in_data_T_1346 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1435 = _fifo_in_data_T_1346 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1446 = _fifo_in_data_T_1346 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1457 = _fifo_in_data_T_1346 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1468 = _fifo_in_data_T_1346 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1479 = _fifo_in_data_T_1346 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1490 = _fifo_in_data_T_1346 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1501 = _fifo_in_data_T_1346 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1512 = _fifo_in_data_T_1346 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1513 = _fifo_in_data_T_1512 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1514 = _fifo_in_data_T_1501 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1513; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1515 = _fifo_in_data_T_1490 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1514; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1516 = _fifo_in_data_T_1479 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1515; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1517 = _fifo_in_data_T_1468 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1516; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1518 = _fifo_in_data_T_1457 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1517; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1519 = _fifo_in_data_T_1446 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1518; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1520 = _fifo_in_data_T_1435 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1519; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1521 = _fifo_in_data_T_1424 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1520; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1522 = _fifo_in_data_T_1413 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1521; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1523 = _fifo_in_data_T_1402 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1522; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1524 = _fifo_in_data_T_1391 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1523; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1525 = _fifo_in_data_T_1380 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1524; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1526 = _fifo_in_data_T_1369 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1525; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1527 = _fifo_in_data_T_1358 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1526; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_7 = _fifo_in_data_T_1347 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1527; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1514 = _fifo_in_data_T_1501 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1512 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1515 = _fifo_in_data_T_1490 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1514; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1516 = _fifo_in_data_T_1479 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1515; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1517 = _fifo_in_data_T_1468 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1516; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1518 = _fifo_in_data_T_1457 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1517; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1519 = _fifo_in_data_T_1446 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1518; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1520 = _fifo_in_data_T_1435 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1519; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1521 = _fifo_in_data_T_1424 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1520; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1522 = _fifo_in_data_T_1413 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1521; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1523 = _fifo_in_data_T_1402 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1522; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1524 = _fifo_in_data_T_1391 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1523; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1525 = _fifo_in_data_T_1380 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1524; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1526 = _fifo_in_data_T_1369 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1525; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1527 = _fifo_in_data_T_1358 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1526; // @[Mux.scala 98:16]
  wire  fifo_in_valid_7 = _fifo_in_data_T_1347 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1527; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1530 = 4'h8 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1534 = _fifo_in_data_T_4 + 5'h8; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1535 = counter <= 4'h8 ? {{1'd0}, _fifo_in_data_T_1530} : _fifo_in_data_T_1534; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1537 = _fifo_in_data_T_1535 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1538 = _fifo_in_data_T_1537 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1549 = _fifo_in_data_T_1537 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1560 = _fifo_in_data_T_1537 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1571 = _fifo_in_data_T_1537 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1582 = _fifo_in_data_T_1537 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1593 = _fifo_in_data_T_1537 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1604 = _fifo_in_data_T_1537 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1615 = _fifo_in_data_T_1537 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1626 = _fifo_in_data_T_1537 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1637 = _fifo_in_data_T_1537 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1648 = _fifo_in_data_T_1537 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1659 = _fifo_in_data_T_1537 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1670 = _fifo_in_data_T_1537 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1681 = _fifo_in_data_T_1537 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1692 = _fifo_in_data_T_1537 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1703 = _fifo_in_data_T_1537 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1704 = _fifo_in_data_T_1703 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1705 = _fifo_in_data_T_1692 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1704; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1706 = _fifo_in_data_T_1681 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1705; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1707 = _fifo_in_data_T_1670 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1706; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1708 = _fifo_in_data_T_1659 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1707; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1709 = _fifo_in_data_T_1648 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1708; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1710 = _fifo_in_data_T_1637 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1709; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1711 = _fifo_in_data_T_1626 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1710; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1712 = _fifo_in_data_T_1615 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1711; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1713 = _fifo_in_data_T_1604 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1712; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1714 = _fifo_in_data_T_1593 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1713; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1715 = _fifo_in_data_T_1582 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1714; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1716 = _fifo_in_data_T_1571 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1715; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1717 = _fifo_in_data_T_1560 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1716; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1718 = _fifo_in_data_T_1549 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1717; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_8 = _fifo_in_data_T_1538 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1718; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1705 = _fifo_in_data_T_1692 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1703 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1706 = _fifo_in_data_T_1681 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1705; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1707 = _fifo_in_data_T_1670 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1706; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1708 = _fifo_in_data_T_1659 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1707; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1709 = _fifo_in_data_T_1648 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1708; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1710 = _fifo_in_data_T_1637 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1709; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1711 = _fifo_in_data_T_1626 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1710; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1712 = _fifo_in_data_T_1615 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1711; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1713 = _fifo_in_data_T_1604 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1712; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1714 = _fifo_in_data_T_1593 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1713; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1715 = _fifo_in_data_T_1582 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1714; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1716 = _fifo_in_data_T_1571 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1715; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1717 = _fifo_in_data_T_1560 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1716; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1718 = _fifo_in_data_T_1549 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1717; // @[Mux.scala 98:16]
  wire  fifo_in_valid_8 = _fifo_in_data_T_1538 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1718; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1721 = 4'h9 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1725 = _fifo_in_data_T_4 + 5'h9; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1726 = counter <= 4'h9 ? {{1'd0}, _fifo_in_data_T_1721} : _fifo_in_data_T_1725; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1728 = _fifo_in_data_T_1726 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1729 = _fifo_in_data_T_1728 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1740 = _fifo_in_data_T_1728 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1751 = _fifo_in_data_T_1728 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1762 = _fifo_in_data_T_1728 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1773 = _fifo_in_data_T_1728 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1784 = _fifo_in_data_T_1728 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1795 = _fifo_in_data_T_1728 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1806 = _fifo_in_data_T_1728 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1817 = _fifo_in_data_T_1728 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1828 = _fifo_in_data_T_1728 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1839 = _fifo_in_data_T_1728 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1850 = _fifo_in_data_T_1728 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1861 = _fifo_in_data_T_1728 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1872 = _fifo_in_data_T_1728 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1883 = _fifo_in_data_T_1728 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1894 = _fifo_in_data_T_1728 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1895 = _fifo_in_data_T_1894 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1896 = _fifo_in_data_T_1883 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1895; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1897 = _fifo_in_data_T_1872 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1896; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1898 = _fifo_in_data_T_1861 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1897; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1899 = _fifo_in_data_T_1850 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1898; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1900 = _fifo_in_data_T_1839 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1899; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1901 = _fifo_in_data_T_1828 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1900; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1902 = _fifo_in_data_T_1817 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1901; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1903 = _fifo_in_data_T_1806 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1902; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1904 = _fifo_in_data_T_1795 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1903; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1905 = _fifo_in_data_T_1784 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1904; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1906 = _fifo_in_data_T_1773 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1905; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1907 = _fifo_in_data_T_1762 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1906; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1908 = _fifo_in_data_T_1751 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1907; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1909 = _fifo_in_data_T_1740 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1908; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_9 = _fifo_in_data_T_1729 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1909; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1896 = _fifo_in_data_T_1883 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1894 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1897 = _fifo_in_data_T_1872 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1896; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1898 = _fifo_in_data_T_1861 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1897; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1899 = _fifo_in_data_T_1850 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1898; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1900 = _fifo_in_data_T_1839 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1899; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1901 = _fifo_in_data_T_1828 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1900; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1902 = _fifo_in_data_T_1817 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1901; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1903 = _fifo_in_data_T_1806 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1902; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1904 = _fifo_in_data_T_1795 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1903; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1905 = _fifo_in_data_T_1784 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1904; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1906 = _fifo_in_data_T_1773 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1905; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1907 = _fifo_in_data_T_1762 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1906; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1908 = _fifo_in_data_T_1751 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1907; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1909 = _fifo_in_data_T_1740 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1908; // @[Mux.scala 98:16]
  wire  fifo_in_valid_9 = _fifo_in_data_T_1729 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1909; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1912 = 4'ha - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1916 = _fifo_in_data_T_4 + 5'ha; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1917 = counter <= 4'ha ? {{1'd0}, _fifo_in_data_T_1912} : _fifo_in_data_T_1916; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1919 = _fifo_in_data_T_1917 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1920 = _fifo_in_data_T_1919 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1931 = _fifo_in_data_T_1919 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1942 = _fifo_in_data_T_1919 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1953 = _fifo_in_data_T_1919 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1964 = _fifo_in_data_T_1919 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1975 = _fifo_in_data_T_1919 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1986 = _fifo_in_data_T_1919 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1997 = _fifo_in_data_T_1919 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2008 = _fifo_in_data_T_1919 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2019 = _fifo_in_data_T_1919 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2030 = _fifo_in_data_T_1919 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2041 = _fifo_in_data_T_1919 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2052 = _fifo_in_data_T_1919 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2063 = _fifo_in_data_T_1919 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2074 = _fifo_in_data_T_1919 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2085 = _fifo_in_data_T_1919 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2086 = _fifo_in_data_T_2085 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2087 = _fifo_in_data_T_2074 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2086; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2088 = _fifo_in_data_T_2063 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2087; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2089 = _fifo_in_data_T_2052 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2088; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2090 = _fifo_in_data_T_2041 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2089; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2091 = _fifo_in_data_T_2030 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2090; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2092 = _fifo_in_data_T_2019 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2091; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2093 = _fifo_in_data_T_2008 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2092; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2094 = _fifo_in_data_T_1997 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2093; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2095 = _fifo_in_data_T_1986 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2094; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2096 = _fifo_in_data_T_1975 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2095; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2097 = _fifo_in_data_T_1964 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2096; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2098 = _fifo_in_data_T_1953 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2097; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2099 = _fifo_in_data_T_1942 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2098; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2100 = _fifo_in_data_T_1931 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2099; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_10 = _fifo_in_data_T_1920 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2100; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2087 = _fifo_in_data_T_2074 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2085 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2088 = _fifo_in_data_T_2063 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2087; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2089 = _fifo_in_data_T_2052 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2088; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2090 = _fifo_in_data_T_2041 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2089; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2091 = _fifo_in_data_T_2030 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2090; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2092 = _fifo_in_data_T_2019 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2091; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2093 = _fifo_in_data_T_2008 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2092; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2094 = _fifo_in_data_T_1997 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2093; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2095 = _fifo_in_data_T_1986 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2094; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2096 = _fifo_in_data_T_1975 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2095; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2097 = _fifo_in_data_T_1964 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2096; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2098 = _fifo_in_data_T_1953 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2097; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2099 = _fifo_in_data_T_1942 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2098; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2100 = _fifo_in_data_T_1931 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2099; // @[Mux.scala 98:16]
  wire  fifo_in_valid_10 = _fifo_in_data_T_1920 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2100; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2103 = 4'hb - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2107 = _fifo_in_data_T_4 + 5'hb; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_2108 = counter <= 4'hb ? {{1'd0}, _fifo_in_data_T_2103} : _fifo_in_data_T_2107; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2110 = _fifo_in_data_T_2108 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2111 = _fifo_in_data_T_2110 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2122 = _fifo_in_data_T_2110 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2133 = _fifo_in_data_T_2110 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2144 = _fifo_in_data_T_2110 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2155 = _fifo_in_data_T_2110 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2166 = _fifo_in_data_T_2110 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2177 = _fifo_in_data_T_2110 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2188 = _fifo_in_data_T_2110 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2199 = _fifo_in_data_T_2110 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2210 = _fifo_in_data_T_2110 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2221 = _fifo_in_data_T_2110 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2232 = _fifo_in_data_T_2110 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2243 = _fifo_in_data_T_2110 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2254 = _fifo_in_data_T_2110 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2265 = _fifo_in_data_T_2110 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2276 = _fifo_in_data_T_2110 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2277 = _fifo_in_data_T_2276 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2278 = _fifo_in_data_T_2265 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2277; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2279 = _fifo_in_data_T_2254 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2278; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2280 = _fifo_in_data_T_2243 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2279; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2281 = _fifo_in_data_T_2232 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2280; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2282 = _fifo_in_data_T_2221 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2281; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2283 = _fifo_in_data_T_2210 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2282; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2284 = _fifo_in_data_T_2199 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2283; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2285 = _fifo_in_data_T_2188 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2284; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2286 = _fifo_in_data_T_2177 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2285; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2287 = _fifo_in_data_T_2166 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2286; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2288 = _fifo_in_data_T_2155 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2287; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2289 = _fifo_in_data_T_2144 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2288; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2290 = _fifo_in_data_T_2133 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2289; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2291 = _fifo_in_data_T_2122 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2290; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_11 = _fifo_in_data_T_2111 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2291; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2278 = _fifo_in_data_T_2265 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2276 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2279 = _fifo_in_data_T_2254 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2278; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2280 = _fifo_in_data_T_2243 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2279; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2281 = _fifo_in_data_T_2232 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2280; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2282 = _fifo_in_data_T_2221 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2281; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2283 = _fifo_in_data_T_2210 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2282; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2284 = _fifo_in_data_T_2199 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2283; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2285 = _fifo_in_data_T_2188 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2284; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2286 = _fifo_in_data_T_2177 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2285; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2287 = _fifo_in_data_T_2166 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2286; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2288 = _fifo_in_data_T_2155 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2287; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2289 = _fifo_in_data_T_2144 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2288; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2290 = _fifo_in_data_T_2133 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2289; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2291 = _fifo_in_data_T_2122 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2290; // @[Mux.scala 98:16]
  wire  fifo_in_valid_11 = _fifo_in_data_T_2111 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2291; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2294 = 4'hc - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2298 = _fifo_in_data_T_4 + 5'hc; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_2299 = counter <= 4'hc ? {{1'd0}, _fifo_in_data_T_2294} : _fifo_in_data_T_2298; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2301 = _fifo_in_data_T_2299 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2302 = _fifo_in_data_T_2301 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2313 = _fifo_in_data_T_2301 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2324 = _fifo_in_data_T_2301 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2335 = _fifo_in_data_T_2301 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2346 = _fifo_in_data_T_2301 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2357 = _fifo_in_data_T_2301 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2368 = _fifo_in_data_T_2301 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2379 = _fifo_in_data_T_2301 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2390 = _fifo_in_data_T_2301 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2401 = _fifo_in_data_T_2301 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2412 = _fifo_in_data_T_2301 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2423 = _fifo_in_data_T_2301 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2434 = _fifo_in_data_T_2301 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2445 = _fifo_in_data_T_2301 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2456 = _fifo_in_data_T_2301 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2467 = _fifo_in_data_T_2301 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2468 = _fifo_in_data_T_2467 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2469 = _fifo_in_data_T_2456 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2468; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2470 = _fifo_in_data_T_2445 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2469; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2471 = _fifo_in_data_T_2434 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2470; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2472 = _fifo_in_data_T_2423 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2471; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2473 = _fifo_in_data_T_2412 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2472; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2474 = _fifo_in_data_T_2401 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2473; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2475 = _fifo_in_data_T_2390 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2474; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2476 = _fifo_in_data_T_2379 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2475; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2477 = _fifo_in_data_T_2368 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2476; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2478 = _fifo_in_data_T_2357 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2477; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2479 = _fifo_in_data_T_2346 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2478; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2480 = _fifo_in_data_T_2335 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2479; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2481 = _fifo_in_data_T_2324 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2480; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2482 = _fifo_in_data_T_2313 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2481; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_12 = _fifo_in_data_T_2302 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2482; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2469 = _fifo_in_data_T_2456 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2467 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2470 = _fifo_in_data_T_2445 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2469; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2471 = _fifo_in_data_T_2434 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2470; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2472 = _fifo_in_data_T_2423 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2471; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2473 = _fifo_in_data_T_2412 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2472; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2474 = _fifo_in_data_T_2401 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2473; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2475 = _fifo_in_data_T_2390 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2474; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2476 = _fifo_in_data_T_2379 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2475; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2477 = _fifo_in_data_T_2368 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2476; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2478 = _fifo_in_data_T_2357 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2477; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2479 = _fifo_in_data_T_2346 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2478; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2480 = _fifo_in_data_T_2335 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2479; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2481 = _fifo_in_data_T_2324 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2480; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2482 = _fifo_in_data_T_2313 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2481; // @[Mux.scala 98:16]
  wire  fifo_in_valid_12 = _fifo_in_data_T_2302 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2482; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2485 = 4'hd - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2489 = _fifo_in_data_T_4 + 5'hd; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_2490 = counter <= 4'hd ? {{1'd0}, _fifo_in_data_T_2485} : _fifo_in_data_T_2489; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2492 = _fifo_in_data_T_2490 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2493 = _fifo_in_data_T_2492 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2504 = _fifo_in_data_T_2492 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2515 = _fifo_in_data_T_2492 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2526 = _fifo_in_data_T_2492 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2537 = _fifo_in_data_T_2492 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2548 = _fifo_in_data_T_2492 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2559 = _fifo_in_data_T_2492 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2570 = _fifo_in_data_T_2492 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2581 = _fifo_in_data_T_2492 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2592 = _fifo_in_data_T_2492 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2603 = _fifo_in_data_T_2492 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2614 = _fifo_in_data_T_2492 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2625 = _fifo_in_data_T_2492 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2636 = _fifo_in_data_T_2492 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2647 = _fifo_in_data_T_2492 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2658 = _fifo_in_data_T_2492 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2659 = _fifo_in_data_T_2658 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2660 = _fifo_in_data_T_2647 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2659; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2661 = _fifo_in_data_T_2636 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2660; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2662 = _fifo_in_data_T_2625 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2661; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2663 = _fifo_in_data_T_2614 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2662; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2664 = _fifo_in_data_T_2603 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2663; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2665 = _fifo_in_data_T_2592 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2664; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2666 = _fifo_in_data_T_2581 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2665; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2667 = _fifo_in_data_T_2570 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2666; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2668 = _fifo_in_data_T_2559 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2667; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2669 = _fifo_in_data_T_2548 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2668; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2670 = _fifo_in_data_T_2537 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2669; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2671 = _fifo_in_data_T_2526 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2670; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2672 = _fifo_in_data_T_2515 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2671; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2673 = _fifo_in_data_T_2504 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2672; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_13 = _fifo_in_data_T_2493 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2673; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2660 = _fifo_in_data_T_2647 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2658 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2661 = _fifo_in_data_T_2636 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2660; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2662 = _fifo_in_data_T_2625 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2661; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2663 = _fifo_in_data_T_2614 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2662; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2664 = _fifo_in_data_T_2603 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2663; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2665 = _fifo_in_data_T_2592 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2664; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2666 = _fifo_in_data_T_2581 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2665; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2667 = _fifo_in_data_T_2570 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2666; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2668 = _fifo_in_data_T_2559 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2667; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2669 = _fifo_in_data_T_2548 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2668; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2670 = _fifo_in_data_T_2537 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2669; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2671 = _fifo_in_data_T_2526 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2670; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2672 = _fifo_in_data_T_2515 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2671; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2673 = _fifo_in_data_T_2504 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2672; // @[Mux.scala 98:16]
  wire  fifo_in_valid_13 = _fifo_in_data_T_2493 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2673; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2676 = 4'he - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2680 = _fifo_in_data_T_4 + 5'he; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_2681 = counter <= 4'he ? {{1'd0}, _fifo_in_data_T_2676} : _fifo_in_data_T_2680; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2683 = _fifo_in_data_T_2681 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2684 = _fifo_in_data_T_2683 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2695 = _fifo_in_data_T_2683 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2706 = _fifo_in_data_T_2683 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2717 = _fifo_in_data_T_2683 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2728 = _fifo_in_data_T_2683 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2739 = _fifo_in_data_T_2683 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2750 = _fifo_in_data_T_2683 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2761 = _fifo_in_data_T_2683 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2772 = _fifo_in_data_T_2683 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2783 = _fifo_in_data_T_2683 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2794 = _fifo_in_data_T_2683 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2805 = _fifo_in_data_T_2683 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2816 = _fifo_in_data_T_2683 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2827 = _fifo_in_data_T_2683 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2838 = _fifo_in_data_T_2683 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2849 = _fifo_in_data_T_2683 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2850 = _fifo_in_data_T_2849 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2851 = _fifo_in_data_T_2838 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2850; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2852 = _fifo_in_data_T_2827 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2851; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2853 = _fifo_in_data_T_2816 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2852; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2854 = _fifo_in_data_T_2805 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2853; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2855 = _fifo_in_data_T_2794 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2854; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2856 = _fifo_in_data_T_2783 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2855; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2857 = _fifo_in_data_T_2772 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2856; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2858 = _fifo_in_data_T_2761 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2857; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2859 = _fifo_in_data_T_2750 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2858; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2860 = _fifo_in_data_T_2739 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2859; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2861 = _fifo_in_data_T_2728 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2860; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2862 = _fifo_in_data_T_2717 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2861; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2863 = _fifo_in_data_T_2706 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2862; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2864 = _fifo_in_data_T_2695 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2863; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_14 = _fifo_in_data_T_2684 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2864; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2851 = _fifo_in_data_T_2838 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2849 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2852 = _fifo_in_data_T_2827 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2851; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2853 = _fifo_in_data_T_2816 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2852; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2854 = _fifo_in_data_T_2805 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2853; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2855 = _fifo_in_data_T_2794 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2854; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2856 = _fifo_in_data_T_2783 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2855; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2857 = _fifo_in_data_T_2772 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2856; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2858 = _fifo_in_data_T_2761 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2857; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2859 = _fifo_in_data_T_2750 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2858; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2860 = _fifo_in_data_T_2739 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2859; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2861 = _fifo_in_data_T_2728 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2860; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2862 = _fifo_in_data_T_2717 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2861; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2863 = _fifo_in_data_T_2706 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2862; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2864 = _fifo_in_data_T_2695 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2863; // @[Mux.scala 98:16]
  wire  fifo_in_valid_14 = _fifo_in_data_T_2684 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2864; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2867 = 4'hf - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2872 = {{1'd0}, _fifo_in_data_T_2867}; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2874 = _fifo_in_data_T_2872 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2875 = _fifo_in_data_T_2874 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2886 = _fifo_in_data_T_2874 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2897 = _fifo_in_data_T_2874 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2908 = _fifo_in_data_T_2874 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2919 = _fifo_in_data_T_2874 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2930 = _fifo_in_data_T_2874 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2941 = _fifo_in_data_T_2874 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2952 = _fifo_in_data_T_2874 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2963 = _fifo_in_data_T_2874 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2974 = _fifo_in_data_T_2874 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2985 = _fifo_in_data_T_2874 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2996 = _fifo_in_data_T_2874 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_3007 = _fifo_in_data_T_2874 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_3018 = _fifo_in_data_T_2874 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_3029 = _fifo_in_data_T_2874 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_3040 = _fifo_in_data_T_2874 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_3041 = _fifo_in_data_T_3040 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3042 = _fifo_in_data_T_3029 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_3041; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3043 = _fifo_in_data_T_3018 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_3042; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3044 = _fifo_in_data_T_3007 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_3043; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3045 = _fifo_in_data_T_2996 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_3044; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3046 = _fifo_in_data_T_2985 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_3045; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3047 = _fifo_in_data_T_2974 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_3046; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3048 = _fifo_in_data_T_2963 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_3047; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3049 = _fifo_in_data_T_2952 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_3048; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3050 = _fifo_in_data_T_2941 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_3049; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3051 = _fifo_in_data_T_2930 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_3050; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3052 = _fifo_in_data_T_2919 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_3051; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3053 = _fifo_in_data_T_2908 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_3052; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3054 = _fifo_in_data_T_2897 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_3053; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3055 = _fifo_in_data_T_2886 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_3054; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_15 = _fifo_in_data_T_2875 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_3055; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3042 = _fifo_in_data_T_3029 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_3040 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3043 = _fifo_in_data_T_3018 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_3042; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3044 = _fifo_in_data_T_3007 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_3043; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3045 = _fifo_in_data_T_2996 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_3044; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3046 = _fifo_in_data_T_2985 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_3045; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3047 = _fifo_in_data_T_2974 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_3046; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3048 = _fifo_in_data_T_2963 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_3047; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3049 = _fifo_in_data_T_2952 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_3048; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3050 = _fifo_in_data_T_2941 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_3049; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3051 = _fifo_in_data_T_2930 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_3050; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3052 = _fifo_in_data_T_2919 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_3051; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3053 = _fifo_in_data_T_2908 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_3052; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3054 = _fifo_in_data_T_2897 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_3053; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3055 = _fifo_in_data_T_2886 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_3054; // @[Mux.scala 98:16]
  wire  fifo_in_valid_15 = _fifo_in_data_T_2875 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_3055; // @[Mux.scala 98:16]
  wire [31:0] collector_data_1 = collector_fifos_1_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_0 = collector_fifos_0_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_3 = collector_fifos_3_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_2 = collector_fifos_2_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_5 = collector_fifos_5_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_4 = collector_fifos_4_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_7 = collector_fifos_7_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_6 = collector_fifos_6_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [255:0] io_out_dout_lo = {collector_data_7,collector_data_6,collector_data_5,collector_data_4,collector_data_3,
    collector_data_2,collector_data_1,collector_data_0}; // @[BFS.scala 877:39]
  wire [31:0] collector_data_9 = collector_fifos_9_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_8 = collector_fifos_8_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_11 = collector_fifos_11_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_10 = collector_fifos_10_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_13 = collector_fifos_13_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_12 = collector_fifos_12_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_15 = collector_fifos_15_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_14 = collector_fifos_14_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [255:0] io_out_dout_hi = {collector_data_15,collector_data_14,collector_data_13,collector_data_12,
    collector_data_11,collector_data_10,collector_data_9,collector_data_8}; // @[BFS.scala 877:39]
  wire [8:0] _io_out_data_count_WIRE = {{4'd0}, collector_fifos_0_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_WIRE_1 = {{4'd0}, collector_fifos_1_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_1 = _io_out_data_count_WIRE + _io_out_data_count_WIRE_1; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_2 = {{4'd0}, collector_fifos_2_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_3 = _io_out_data_count_T_1 + _io_out_data_count_WIRE_2; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_3 = {{4'd0}, collector_fifos_3_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_5 = _io_out_data_count_T_3 + _io_out_data_count_WIRE_3; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_4 = {{4'd0}, collector_fifos_4_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_7 = _io_out_data_count_T_5 + _io_out_data_count_WIRE_4; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_5 = {{4'd0}, collector_fifos_5_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_9 = _io_out_data_count_T_7 + _io_out_data_count_WIRE_5; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_6 = {{4'd0}, collector_fifos_6_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_11 = _io_out_data_count_T_9 + _io_out_data_count_WIRE_6; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_7 = {{4'd0}, collector_fifos_7_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_13 = _io_out_data_count_T_11 + _io_out_data_count_WIRE_7; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_8 = {{4'd0}, collector_fifos_8_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_15 = _io_out_data_count_T_13 + _io_out_data_count_WIRE_8; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_9 = {{4'd0}, collector_fifos_9_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_17 = _io_out_data_count_T_15 + _io_out_data_count_WIRE_9; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_10 = {{4'd0}, collector_fifos_10_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_19 = _io_out_data_count_T_17 + _io_out_data_count_WIRE_10; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_11 = {{4'd0}, collector_fifos_11_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_21 = _io_out_data_count_T_19 + _io_out_data_count_WIRE_11; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_12 = {{4'd0}, collector_fifos_12_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_23 = _io_out_data_count_T_21 + _io_out_data_count_WIRE_12; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_13 = {{4'd0}, collector_fifos_13_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_25 = _io_out_data_count_T_23 + _io_out_data_count_WIRE_13; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_14 = {{4'd0}, collector_fifos_14_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_27 = _io_out_data_count_T_25 + _io_out_data_count_WIRE_14; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_15 = {{4'd0}, collector_fifos_15_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  collector_fifo_0 collector_fifos_0 ( // @[BFS.scala 826:16]
    .full(collector_fifos_0_full),
    .din(collector_fifos_0_din),
    .wr_en(collector_fifos_0_wr_en),
    .empty(collector_fifos_0_empty),
    .dout(collector_fifos_0_dout),
    .rd_en(collector_fifos_0_rd_en),
    .data_count(collector_fifos_0_data_count),
    .clk(collector_fifos_0_clk),
    .srst(collector_fifos_0_srst),
    .valid(collector_fifos_0_valid)
  );
  collector_fifo_0 collector_fifos_1 ( // @[BFS.scala 826:16]
    .full(collector_fifos_1_full),
    .din(collector_fifos_1_din),
    .wr_en(collector_fifos_1_wr_en),
    .empty(collector_fifos_1_empty),
    .dout(collector_fifos_1_dout),
    .rd_en(collector_fifos_1_rd_en),
    .data_count(collector_fifos_1_data_count),
    .clk(collector_fifos_1_clk),
    .srst(collector_fifos_1_srst),
    .valid(collector_fifos_1_valid)
  );
  collector_fifo_0 collector_fifos_2 ( // @[BFS.scala 826:16]
    .full(collector_fifos_2_full),
    .din(collector_fifos_2_din),
    .wr_en(collector_fifos_2_wr_en),
    .empty(collector_fifos_2_empty),
    .dout(collector_fifos_2_dout),
    .rd_en(collector_fifos_2_rd_en),
    .data_count(collector_fifos_2_data_count),
    .clk(collector_fifos_2_clk),
    .srst(collector_fifos_2_srst),
    .valid(collector_fifos_2_valid)
  );
  collector_fifo_0 collector_fifos_3 ( // @[BFS.scala 826:16]
    .full(collector_fifos_3_full),
    .din(collector_fifos_3_din),
    .wr_en(collector_fifos_3_wr_en),
    .empty(collector_fifos_3_empty),
    .dout(collector_fifos_3_dout),
    .rd_en(collector_fifos_3_rd_en),
    .data_count(collector_fifos_3_data_count),
    .clk(collector_fifos_3_clk),
    .srst(collector_fifos_3_srst),
    .valid(collector_fifos_3_valid)
  );
  collector_fifo_0 collector_fifos_4 ( // @[BFS.scala 826:16]
    .full(collector_fifos_4_full),
    .din(collector_fifos_4_din),
    .wr_en(collector_fifos_4_wr_en),
    .empty(collector_fifos_4_empty),
    .dout(collector_fifos_4_dout),
    .rd_en(collector_fifos_4_rd_en),
    .data_count(collector_fifos_4_data_count),
    .clk(collector_fifos_4_clk),
    .srst(collector_fifos_4_srst),
    .valid(collector_fifos_4_valid)
  );
  collector_fifo_0 collector_fifos_5 ( // @[BFS.scala 826:16]
    .full(collector_fifos_5_full),
    .din(collector_fifos_5_din),
    .wr_en(collector_fifos_5_wr_en),
    .empty(collector_fifos_5_empty),
    .dout(collector_fifos_5_dout),
    .rd_en(collector_fifos_5_rd_en),
    .data_count(collector_fifos_5_data_count),
    .clk(collector_fifos_5_clk),
    .srst(collector_fifos_5_srst),
    .valid(collector_fifos_5_valid)
  );
  collector_fifo_0 collector_fifos_6 ( // @[BFS.scala 826:16]
    .full(collector_fifos_6_full),
    .din(collector_fifos_6_din),
    .wr_en(collector_fifos_6_wr_en),
    .empty(collector_fifos_6_empty),
    .dout(collector_fifos_6_dout),
    .rd_en(collector_fifos_6_rd_en),
    .data_count(collector_fifos_6_data_count),
    .clk(collector_fifos_6_clk),
    .srst(collector_fifos_6_srst),
    .valid(collector_fifos_6_valid)
  );
  collector_fifo_0 collector_fifos_7 ( // @[BFS.scala 826:16]
    .full(collector_fifos_7_full),
    .din(collector_fifos_7_din),
    .wr_en(collector_fifos_7_wr_en),
    .empty(collector_fifos_7_empty),
    .dout(collector_fifos_7_dout),
    .rd_en(collector_fifos_7_rd_en),
    .data_count(collector_fifos_7_data_count),
    .clk(collector_fifos_7_clk),
    .srst(collector_fifos_7_srst),
    .valid(collector_fifos_7_valid)
  );
  collector_fifo_0 collector_fifos_8 ( // @[BFS.scala 826:16]
    .full(collector_fifos_8_full),
    .din(collector_fifos_8_din),
    .wr_en(collector_fifos_8_wr_en),
    .empty(collector_fifos_8_empty),
    .dout(collector_fifos_8_dout),
    .rd_en(collector_fifos_8_rd_en),
    .data_count(collector_fifos_8_data_count),
    .clk(collector_fifos_8_clk),
    .srst(collector_fifos_8_srst),
    .valid(collector_fifos_8_valid)
  );
  collector_fifo_0 collector_fifos_9 ( // @[BFS.scala 826:16]
    .full(collector_fifos_9_full),
    .din(collector_fifos_9_din),
    .wr_en(collector_fifos_9_wr_en),
    .empty(collector_fifos_9_empty),
    .dout(collector_fifos_9_dout),
    .rd_en(collector_fifos_9_rd_en),
    .data_count(collector_fifos_9_data_count),
    .clk(collector_fifos_9_clk),
    .srst(collector_fifos_9_srst),
    .valid(collector_fifos_9_valid)
  );
  collector_fifo_0 collector_fifos_10 ( // @[BFS.scala 826:16]
    .full(collector_fifos_10_full),
    .din(collector_fifos_10_din),
    .wr_en(collector_fifos_10_wr_en),
    .empty(collector_fifos_10_empty),
    .dout(collector_fifos_10_dout),
    .rd_en(collector_fifos_10_rd_en),
    .data_count(collector_fifos_10_data_count),
    .clk(collector_fifos_10_clk),
    .srst(collector_fifos_10_srst),
    .valid(collector_fifos_10_valid)
  );
  collector_fifo_0 collector_fifos_11 ( // @[BFS.scala 826:16]
    .full(collector_fifos_11_full),
    .din(collector_fifos_11_din),
    .wr_en(collector_fifos_11_wr_en),
    .empty(collector_fifos_11_empty),
    .dout(collector_fifos_11_dout),
    .rd_en(collector_fifos_11_rd_en),
    .data_count(collector_fifos_11_data_count),
    .clk(collector_fifos_11_clk),
    .srst(collector_fifos_11_srst),
    .valid(collector_fifos_11_valid)
  );
  collector_fifo_0 collector_fifos_12 ( // @[BFS.scala 826:16]
    .full(collector_fifos_12_full),
    .din(collector_fifos_12_din),
    .wr_en(collector_fifos_12_wr_en),
    .empty(collector_fifos_12_empty),
    .dout(collector_fifos_12_dout),
    .rd_en(collector_fifos_12_rd_en),
    .data_count(collector_fifos_12_data_count),
    .clk(collector_fifos_12_clk),
    .srst(collector_fifos_12_srst),
    .valid(collector_fifos_12_valid)
  );
  collector_fifo_0 collector_fifos_13 ( // @[BFS.scala 826:16]
    .full(collector_fifos_13_full),
    .din(collector_fifos_13_din),
    .wr_en(collector_fifos_13_wr_en),
    .empty(collector_fifos_13_empty),
    .dout(collector_fifos_13_dout),
    .rd_en(collector_fifos_13_rd_en),
    .data_count(collector_fifos_13_data_count),
    .clk(collector_fifos_13_clk),
    .srst(collector_fifos_13_srst),
    .valid(collector_fifos_13_valid)
  );
  collector_fifo_0 collector_fifos_14 ( // @[BFS.scala 826:16]
    .full(collector_fifos_14_full),
    .din(collector_fifos_14_din),
    .wr_en(collector_fifos_14_wr_en),
    .empty(collector_fifos_14_empty),
    .dout(collector_fifos_14_dout),
    .rd_en(collector_fifos_14_rd_en),
    .data_count(collector_fifos_14_data_count),
    .clk(collector_fifos_14_clk),
    .srst(collector_fifos_14_srst),
    .valid(collector_fifos_14_valid)
  );
  collector_fifo_0 collector_fifos_15 ( // @[BFS.scala 826:16]
    .full(collector_fifos_15_full),
    .din(collector_fifos_15_din),
    .wr_en(collector_fifos_15_wr_en),
    .empty(collector_fifos_15_empty),
    .dout(collector_fifos_15_dout),
    .rd_en(collector_fifos_15_rd_en),
    .data_count(collector_fifos_15_data_count),
    .clk(collector_fifos_15_clk),
    .srst(collector_fifos_15_srst),
    .valid(collector_fifos_15_valid)
  );
  pipeline in_pipeline_0 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_0_clock),
    .reset(in_pipeline_0_reset),
    .io_dout_ready(in_pipeline_0_io_dout_ready),
    .io_dout_valid(in_pipeline_0_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_0_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_0_io_din_ready),
    .io_din_valid(in_pipeline_0_io_din_valid),
    .io_din_bits_tdata(in_pipeline_0_io_din_bits_tdata)
  );
  pipeline in_pipeline_1 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_1_clock),
    .reset(in_pipeline_1_reset),
    .io_dout_ready(in_pipeline_1_io_dout_ready),
    .io_dout_valid(in_pipeline_1_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_1_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_1_io_din_ready),
    .io_din_valid(in_pipeline_1_io_din_valid),
    .io_din_bits_tdata(in_pipeline_1_io_din_bits_tdata)
  );
  pipeline in_pipeline_2 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_2_clock),
    .reset(in_pipeline_2_reset),
    .io_dout_ready(in_pipeline_2_io_dout_ready),
    .io_dout_valid(in_pipeline_2_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_2_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_2_io_din_ready),
    .io_din_valid(in_pipeline_2_io_din_valid),
    .io_din_bits_tdata(in_pipeline_2_io_din_bits_tdata)
  );
  pipeline in_pipeline_3 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_3_clock),
    .reset(in_pipeline_3_reset),
    .io_dout_ready(in_pipeline_3_io_dout_ready),
    .io_dout_valid(in_pipeline_3_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_3_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_3_io_din_ready),
    .io_din_valid(in_pipeline_3_io_din_valid),
    .io_din_bits_tdata(in_pipeline_3_io_din_bits_tdata)
  );
  pipeline in_pipeline_4 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_4_clock),
    .reset(in_pipeline_4_reset),
    .io_dout_ready(in_pipeline_4_io_dout_ready),
    .io_dout_valid(in_pipeline_4_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_4_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_4_io_din_ready),
    .io_din_valid(in_pipeline_4_io_din_valid),
    .io_din_bits_tdata(in_pipeline_4_io_din_bits_tdata)
  );
  pipeline in_pipeline_5 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_5_clock),
    .reset(in_pipeline_5_reset),
    .io_dout_ready(in_pipeline_5_io_dout_ready),
    .io_dout_valid(in_pipeline_5_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_5_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_5_io_din_ready),
    .io_din_valid(in_pipeline_5_io_din_valid),
    .io_din_bits_tdata(in_pipeline_5_io_din_bits_tdata)
  );
  pipeline in_pipeline_6 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_6_clock),
    .reset(in_pipeline_6_reset),
    .io_dout_ready(in_pipeline_6_io_dout_ready),
    .io_dout_valid(in_pipeline_6_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_6_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_6_io_din_ready),
    .io_din_valid(in_pipeline_6_io_din_valid),
    .io_din_bits_tdata(in_pipeline_6_io_din_bits_tdata)
  );
  pipeline in_pipeline_7 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_7_clock),
    .reset(in_pipeline_7_reset),
    .io_dout_ready(in_pipeline_7_io_dout_ready),
    .io_dout_valid(in_pipeline_7_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_7_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_7_io_din_ready),
    .io_din_valid(in_pipeline_7_io_din_valid),
    .io_din_bits_tdata(in_pipeline_7_io_din_bits_tdata)
  );
  pipeline in_pipeline_8 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_8_clock),
    .reset(in_pipeline_8_reset),
    .io_dout_ready(in_pipeline_8_io_dout_ready),
    .io_dout_valid(in_pipeline_8_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_8_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_8_io_din_ready),
    .io_din_valid(in_pipeline_8_io_din_valid),
    .io_din_bits_tdata(in_pipeline_8_io_din_bits_tdata)
  );
  pipeline in_pipeline_9 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_9_clock),
    .reset(in_pipeline_9_reset),
    .io_dout_ready(in_pipeline_9_io_dout_ready),
    .io_dout_valid(in_pipeline_9_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_9_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_9_io_din_ready),
    .io_din_valid(in_pipeline_9_io_din_valid),
    .io_din_bits_tdata(in_pipeline_9_io_din_bits_tdata)
  );
  pipeline in_pipeline_10 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_10_clock),
    .reset(in_pipeline_10_reset),
    .io_dout_ready(in_pipeline_10_io_dout_ready),
    .io_dout_valid(in_pipeline_10_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_10_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_10_io_din_ready),
    .io_din_valid(in_pipeline_10_io_din_valid),
    .io_din_bits_tdata(in_pipeline_10_io_din_bits_tdata)
  );
  pipeline in_pipeline_11 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_11_clock),
    .reset(in_pipeline_11_reset),
    .io_dout_ready(in_pipeline_11_io_dout_ready),
    .io_dout_valid(in_pipeline_11_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_11_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_11_io_din_ready),
    .io_din_valid(in_pipeline_11_io_din_valid),
    .io_din_bits_tdata(in_pipeline_11_io_din_bits_tdata)
  );
  pipeline in_pipeline_12 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_12_clock),
    .reset(in_pipeline_12_reset),
    .io_dout_ready(in_pipeline_12_io_dout_ready),
    .io_dout_valid(in_pipeline_12_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_12_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_12_io_din_ready),
    .io_din_valid(in_pipeline_12_io_din_valid),
    .io_din_bits_tdata(in_pipeline_12_io_din_bits_tdata)
  );
  pipeline in_pipeline_13 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_13_clock),
    .reset(in_pipeline_13_reset),
    .io_dout_ready(in_pipeline_13_io_dout_ready),
    .io_dout_valid(in_pipeline_13_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_13_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_13_io_din_ready),
    .io_din_valid(in_pipeline_13_io_din_valid),
    .io_din_bits_tdata(in_pipeline_13_io_din_bits_tdata)
  );
  pipeline in_pipeline_14 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_14_clock),
    .reset(in_pipeline_14_reset),
    .io_dout_ready(in_pipeline_14_io_dout_ready),
    .io_dout_valid(in_pipeline_14_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_14_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_14_io_din_ready),
    .io_din_valid(in_pipeline_14_io_din_valid),
    .io_din_bits_tdata(in_pipeline_14_io_din_bits_tdata)
  );
  pipeline in_pipeline_15 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_15_clock),
    .reset(in_pipeline_15_reset),
    .io_dout_ready(in_pipeline_15_io_dout_ready),
    .io_dout_valid(in_pipeline_15_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_15_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_15_io_din_ready),
    .io_din_valid(in_pipeline_15_io_din_valid),
    .io_din_bits_tdata(in_pipeline_15_io_din_bits_tdata)
  );
  assign io_in_0_ready = in_pipeline_0_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_1_ready = in_pipeline_1_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_2_ready = in_pipeline_2_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_3_ready = in_pipeline_3_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_4_ready = in_pipeline_4_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_5_ready = in_pipeline_5_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_6_ready = in_pipeline_6_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_7_ready = in_pipeline_7_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_8_ready = in_pipeline_8_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_9_ready = in_pipeline_9_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_10_ready = in_pipeline_10_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_11_ready = in_pipeline_11_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_12_ready = in_pipeline_12_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_13_ready = in_pipeline_13_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_14_ready = in_pipeline_14_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_15_ready = in_pipeline_15_io_din_ready; // @[BFS.scala 836:16]
  assign io_out_full = ~fifos_ready; // @[BFS.scala 879:18]
  assign io_out_dout = {io_out_dout_hi,io_out_dout_lo}; // @[BFS.scala 877:39]
  assign io_out_data_count = _io_out_data_count_T_27 + _io_out_data_count_WIRE_15; // @[BFS.scala 878:134]
  assign io_out_valid = collector_fifos_0_valid | collector_fifos_1_valid | collector_fifos_2_valid |
    collector_fifos_3_valid | collector_fifos_4_valid | collector_fifos_5_valid | collector_fifos_6_valid |
    collector_fifos_7_valid | collector_fifos_8_valid | collector_fifos_9_valid | collector_fifos_10_valid |
    collector_fifos_11_valid | collector_fifos_12_valid | collector_fifos_13_valid | collector_fifos_14_valid |
    collector_fifos_15_valid; // @[BFS.scala 876:80]
  assign collector_fifos_0_din = io_is_current_tier ? io_out_din[31:0] : fifo_in_data; // @[BFS.scala 867:22]
  assign collector_fifos_0_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid; // @[BFS.scala 868:24]
  assign collector_fifos_0_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_0_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_0_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_1_din = io_is_current_tier ? io_out_din[63:32] : fifo_in_data_1; // @[BFS.scala 867:22]
  assign collector_fifos_1_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_1; // @[BFS.scala 868:24]
  assign collector_fifos_1_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_1_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_1_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_2_din = io_is_current_tier ? io_out_din[95:64] : fifo_in_data_2; // @[BFS.scala 867:22]
  assign collector_fifos_2_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_2; // @[BFS.scala 868:24]
  assign collector_fifos_2_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_2_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_2_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_3_din = io_is_current_tier ? io_out_din[127:96] : fifo_in_data_3; // @[BFS.scala 867:22]
  assign collector_fifos_3_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_3; // @[BFS.scala 868:24]
  assign collector_fifos_3_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_3_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_3_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_4_din = io_is_current_tier ? io_out_din[159:128] : fifo_in_data_4; // @[BFS.scala 867:22]
  assign collector_fifos_4_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_4; // @[BFS.scala 868:24]
  assign collector_fifos_4_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_4_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_4_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_5_din = io_is_current_tier ? io_out_din[191:160] : fifo_in_data_5; // @[BFS.scala 867:22]
  assign collector_fifos_5_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_5; // @[BFS.scala 868:24]
  assign collector_fifos_5_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_5_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_5_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_6_din = io_is_current_tier ? io_out_din[223:192] : fifo_in_data_6; // @[BFS.scala 867:22]
  assign collector_fifos_6_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_6; // @[BFS.scala 868:24]
  assign collector_fifos_6_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_6_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_6_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_7_din = io_is_current_tier ? io_out_din[255:224] : fifo_in_data_7; // @[BFS.scala 867:22]
  assign collector_fifos_7_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_7; // @[BFS.scala 868:24]
  assign collector_fifos_7_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_7_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_7_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_8_din = io_is_current_tier ? io_out_din[287:256] : fifo_in_data_8; // @[BFS.scala 867:22]
  assign collector_fifos_8_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_8; // @[BFS.scala 868:24]
  assign collector_fifos_8_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_8_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_8_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_9_din = io_is_current_tier ? io_out_din[319:288] : fifo_in_data_9; // @[BFS.scala 867:22]
  assign collector_fifos_9_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_9; // @[BFS.scala 868:24]
  assign collector_fifos_9_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_9_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_9_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_10_din = io_is_current_tier ? io_out_din[351:320] : fifo_in_data_10; // @[BFS.scala 867:22]
  assign collector_fifos_10_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_10; // @[BFS.scala 868:24]
  assign collector_fifos_10_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_10_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_10_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_11_din = io_is_current_tier ? io_out_din[383:352] : fifo_in_data_11; // @[BFS.scala 867:22]
  assign collector_fifos_11_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_11; // @[BFS.scala 868:24]
  assign collector_fifos_11_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_11_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_11_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_12_din = io_is_current_tier ? io_out_din[415:384] : fifo_in_data_12; // @[BFS.scala 867:22]
  assign collector_fifos_12_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_12; // @[BFS.scala 868:24]
  assign collector_fifos_12_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_12_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_12_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_13_din = io_is_current_tier ? io_out_din[447:416] : fifo_in_data_13; // @[BFS.scala 867:22]
  assign collector_fifos_13_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_13; // @[BFS.scala 868:24]
  assign collector_fifos_13_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_13_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_13_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_14_din = io_is_current_tier ? io_out_din[479:448] : fifo_in_data_14; // @[BFS.scala 867:22]
  assign collector_fifos_14_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_14; // @[BFS.scala 868:24]
  assign collector_fifos_14_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_14_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_14_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_15_din = io_is_current_tier ? io_out_din[511:480] : fifo_in_data_15; // @[BFS.scala 867:22]
  assign collector_fifos_15_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_15; // @[BFS.scala 868:24]
  assign collector_fifos_15_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_15_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_15_srst = reset; // @[BFS.scala 871:32]
  assign in_pipeline_0_clock = clock;
  assign in_pipeline_0_reset = reset;
  assign in_pipeline_0_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_0_io_din_valid = io_in_0_valid; // @[BFS.scala 836:16]
  assign in_pipeline_0_io_din_bits_tdata = io_in_0_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_1_clock = clock;
  assign in_pipeline_1_reset = reset;
  assign in_pipeline_1_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_1_io_din_valid = io_in_1_valid; // @[BFS.scala 836:16]
  assign in_pipeline_1_io_din_bits_tdata = io_in_1_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_2_clock = clock;
  assign in_pipeline_2_reset = reset;
  assign in_pipeline_2_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_2_io_din_valid = io_in_2_valid; // @[BFS.scala 836:16]
  assign in_pipeline_2_io_din_bits_tdata = io_in_2_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_3_clock = clock;
  assign in_pipeline_3_reset = reset;
  assign in_pipeline_3_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_3_io_din_valid = io_in_3_valid; // @[BFS.scala 836:16]
  assign in_pipeline_3_io_din_bits_tdata = io_in_3_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_4_clock = clock;
  assign in_pipeline_4_reset = reset;
  assign in_pipeline_4_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_4_io_din_valid = io_in_4_valid; // @[BFS.scala 836:16]
  assign in_pipeline_4_io_din_bits_tdata = io_in_4_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_5_clock = clock;
  assign in_pipeline_5_reset = reset;
  assign in_pipeline_5_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_5_io_din_valid = io_in_5_valid; // @[BFS.scala 836:16]
  assign in_pipeline_5_io_din_bits_tdata = io_in_5_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_6_clock = clock;
  assign in_pipeline_6_reset = reset;
  assign in_pipeline_6_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_6_io_din_valid = io_in_6_valid; // @[BFS.scala 836:16]
  assign in_pipeline_6_io_din_bits_tdata = io_in_6_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_7_clock = clock;
  assign in_pipeline_7_reset = reset;
  assign in_pipeline_7_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_7_io_din_valid = io_in_7_valid; // @[BFS.scala 836:16]
  assign in_pipeline_7_io_din_bits_tdata = io_in_7_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_8_clock = clock;
  assign in_pipeline_8_reset = reset;
  assign in_pipeline_8_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_8_io_din_valid = io_in_8_valid; // @[BFS.scala 836:16]
  assign in_pipeline_8_io_din_bits_tdata = io_in_8_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_9_clock = clock;
  assign in_pipeline_9_reset = reset;
  assign in_pipeline_9_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_9_io_din_valid = io_in_9_valid; // @[BFS.scala 836:16]
  assign in_pipeline_9_io_din_bits_tdata = io_in_9_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_10_clock = clock;
  assign in_pipeline_10_reset = reset;
  assign in_pipeline_10_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_10_io_din_valid = io_in_10_valid; // @[BFS.scala 836:16]
  assign in_pipeline_10_io_din_bits_tdata = io_in_10_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_11_clock = clock;
  assign in_pipeline_11_reset = reset;
  assign in_pipeline_11_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_11_io_din_valid = io_in_11_valid; // @[BFS.scala 836:16]
  assign in_pipeline_11_io_din_bits_tdata = io_in_11_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_12_clock = clock;
  assign in_pipeline_12_reset = reset;
  assign in_pipeline_12_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_12_io_din_valid = io_in_12_valid; // @[BFS.scala 836:16]
  assign in_pipeline_12_io_din_bits_tdata = io_in_12_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_13_clock = clock;
  assign in_pipeline_13_reset = reset;
  assign in_pipeline_13_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_13_io_din_valid = io_in_13_valid; // @[BFS.scala 836:16]
  assign in_pipeline_13_io_din_bits_tdata = io_in_13_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_14_clock = clock;
  assign in_pipeline_14_reset = reset;
  assign in_pipeline_14_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_14_io_din_valid = io_in_14_valid; // @[BFS.scala 836:16]
  assign in_pipeline_14_io_din_bits_tdata = io_in_14_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_15_clock = clock;
  assign in_pipeline_15_reset = reset;
  assign in_pipeline_15_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_15_io_din_valid = io_in_15_valid; // @[BFS.scala 836:16]
  assign in_pipeline_15_io_din_bits_tdata = io_in_15_bits_tdata; // @[BFS.scala 836:16]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 829:24]
      counter <= 4'h0; // @[BFS.scala 829:24]
    end else begin
      counter <= _GEN_1[3:0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multi_port_mc(
  input          clock,
  input          reset,
  input          io_cacheable_out_ready,
  output         io_cacheable_out_valid,
  output [511:0] io_cacheable_out_bits_tdata,
  output [15:0]  io_cacheable_out_bits_tkeep,
  output         io_cacheable_in_0_ready,
  input          io_cacheable_in_0_valid,
  input  [31:0]  io_cacheable_in_0_bits_tdata,
  output         io_cacheable_in_1_ready,
  input          io_cacheable_in_1_valid,
  input  [31:0]  io_cacheable_in_1_bits_tdata,
  output         io_cacheable_in_2_ready,
  input          io_cacheable_in_2_valid,
  input  [31:0]  io_cacheable_in_2_bits_tdata,
  output         io_cacheable_in_3_ready,
  input          io_cacheable_in_3_valid,
  input  [31:0]  io_cacheable_in_3_bits_tdata,
  output         io_cacheable_in_4_ready,
  input          io_cacheable_in_4_valid,
  input  [31:0]  io_cacheable_in_4_bits_tdata,
  output         io_cacheable_in_5_ready,
  input          io_cacheable_in_5_valid,
  input  [31:0]  io_cacheable_in_5_bits_tdata,
  output         io_cacheable_in_6_ready,
  input          io_cacheable_in_6_valid,
  input  [31:0]  io_cacheable_in_6_bits_tdata,
  output         io_cacheable_in_7_ready,
  input          io_cacheable_in_7_valid,
  input  [31:0]  io_cacheable_in_7_bits_tdata,
  output         io_cacheable_in_8_ready,
  input          io_cacheable_in_8_valid,
  input  [31:0]  io_cacheable_in_8_bits_tdata,
  output         io_cacheable_in_9_ready,
  input          io_cacheable_in_9_valid,
  input  [31:0]  io_cacheable_in_9_bits_tdata,
  output         io_cacheable_in_10_ready,
  input          io_cacheable_in_10_valid,
  input  [31:0]  io_cacheable_in_10_bits_tdata,
  output         io_cacheable_in_11_ready,
  input          io_cacheable_in_11_valid,
  input  [31:0]  io_cacheable_in_11_bits_tdata,
  output         io_cacheable_in_12_ready,
  input          io_cacheable_in_12_valid,
  input  [31:0]  io_cacheable_in_12_bits_tdata,
  output         io_cacheable_in_13_ready,
  input          io_cacheable_in_13_valid,
  input  [31:0]  io_cacheable_in_13_bits_tdata,
  output         io_cacheable_in_14_ready,
  input          io_cacheable_in_14_valid,
  input  [31:0]  io_cacheable_in_14_bits_tdata,
  output         io_cacheable_in_15_ready,
  input          io_cacheable_in_15_valid,
  input  [31:0]  io_cacheable_in_15_bits_tdata,
  output         io_non_cacheable_in_aw_ready,
  input          io_non_cacheable_in_aw_valid,
  input  [63:0]  io_non_cacheable_in_aw_bits_awaddr,
  input  [6:0]   io_non_cacheable_in_aw_bits_awid,
  output         io_non_cacheable_in_w_ready,
  input          io_non_cacheable_in_w_valid,
  input  [511:0] io_non_cacheable_in_w_bits_wdata,
  input  [63:0]  io_non_cacheable_in_w_bits_wstrb,
  input          io_ddr_out_0_aw_ready,
  output         io_ddr_out_0_aw_valid,
  output [63:0]  io_ddr_out_0_aw_bits_awaddr,
  input          io_ddr_out_0_ar_ready,
  output         io_ddr_out_0_ar_valid,
  output [63:0]  io_ddr_out_0_ar_bits_araddr,
  input          io_ddr_out_0_w_ready,
  output         io_ddr_out_0_w_valid,
  output [511:0] io_ddr_out_0_w_bits_wdata,
  output         io_ddr_out_0_w_bits_wlast,
  input          io_ddr_out_0_r_valid,
  input  [511:0] io_ddr_out_0_r_bits_rdata,
  input          io_ddr_out_0_r_bits_rlast,
  input          io_ddr_out_1_aw_ready,
  output         io_ddr_out_1_aw_valid,
  output [63:0]  io_ddr_out_1_aw_bits_awaddr,
  output [6:0]   io_ddr_out_1_aw_bits_awid,
  input          io_ddr_out_1_w_ready,
  output         io_ddr_out_1_w_valid,
  output [511:0] io_ddr_out_1_w_bits_wdata,
  output [63:0]  io_ddr_out_1_w_bits_wstrb,
  input  [63:0]  io_tiers_base_addr_0,
  input  [63:0]  io_tiers_base_addr_1,
  output [31:0]  io_unvisited_size,
  input          io_start,
  input          io_signal,
  input          io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  tier_fifo_0_clock; // @[BFS.scala 903:46]
  wire  tier_fifo_0_reset; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_0_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_0_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_0_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_1_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_1_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_1_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_2_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_2_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_2_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_3_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_3_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_3_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_4_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_4_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_4_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_5_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_5_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_5_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_6_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_6_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_6_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_7_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_7_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_7_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_8_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_8_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_8_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_9_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_9_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_9_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_10_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_10_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_10_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_11_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_11_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_11_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_12_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_12_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_12_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_13_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_13_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_13_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_14_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_14_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_14_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_15_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_15_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_15_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_out_full; // @[BFS.scala 903:46]
  wire [511:0] tier_fifo_0_io_out_din; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_out_wr_en; // @[BFS.scala 903:46]
  wire [511:0] tier_fifo_0_io_out_dout; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_out_rd_en; // @[BFS.scala 903:46]
  wire [8:0] tier_fifo_0_io_out_data_count; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_out_valid; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_flush; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_is_current_tier; // @[BFS.scala 903:46]
  wire  tier_fifo_1_clock; // @[BFS.scala 903:46]
  wire  tier_fifo_1_reset; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_0_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_0_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_0_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_1_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_1_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_1_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_2_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_2_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_2_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_3_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_3_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_3_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_4_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_4_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_4_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_5_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_5_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_5_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_6_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_6_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_6_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_7_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_7_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_7_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_8_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_8_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_8_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_9_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_9_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_9_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_10_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_10_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_10_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_11_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_11_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_11_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_12_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_12_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_12_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_13_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_13_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_13_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_14_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_14_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_14_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_15_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_15_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_15_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_out_full; // @[BFS.scala 903:46]
  wire [511:0] tier_fifo_1_io_out_din; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_out_wr_en; // @[BFS.scala 903:46]
  wire [511:0] tier_fifo_1_io_out_dout; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_out_rd_en; // @[BFS.scala 903:46]
  wire [8:0] tier_fifo_1_io_out_data_count; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_out_valid; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_flush; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_is_current_tier; // @[BFS.scala 903:46]
  reg [31:0] tier_counter_0; // @[BFS.scala 904:29]
  reg [31:0] tier_counter_1; // @[BFS.scala 904:29]
  reg [4:0] status; // @[BFS.scala 922:23]
  reg [4:0] tier_status_0; // @[BFS.scala 923:28]
  reg [4:0] tier_status_1; // @[BFS.scala 923:28]
  wire  _T_1 = io_start & status == 5'h0; // @[BFS.scala 925:17]
  wire  _T_2 = status == 5'h2; // @[BFS.scala 927:21]
  wire  _T_5 = status == 5'h5; // @[BFS.scala 929:21]
  wire  _T_8 = status == 5'h7; // @[BFS.scala 931:34]
  wire [4:0] _GEN_0 = tier_status_1 != 5'h0 ? 5'h12 : 5'h1; // @[BFS.scala 932:39 BFS.scala 933:14 BFS.scala 935:14]
  wire  _T_11 = status == 5'h1; // @[BFS.scala 937:21]
  wire  _T_14 = status == 5'h6; // @[BFS.scala 939:21]
  wire  _T_17 = status == 5'h8; // @[BFS.scala 941:34]
  wire [4:0] _GEN_1 = tier_status_0 != 5'h0 ? 5'h11 : 5'h2; // @[BFS.scala 942:38 BFS.scala 943:14 BFS.scala 945:14]
  wire  _T_20 = status == 5'h11; // @[BFS.scala 947:21]
  wire  _T_21 = tier_status_0 == 5'h0; // @[BFS.scala 947:60]
  wire  _T_23 = status == 5'h12; // @[BFS.scala 949:21]
  wire  _T_24 = tier_status_1 == 5'h0; // @[BFS.scala 949:60]
  wire [4:0] _GEN_2 = io_end ? 5'h0 : status; // @[BFS.scala 951:21 BFS.scala 952:12 BFS.scala 922:23]
  wire [4:0] _GEN_3 = status == 5'h12 & tier_status_1 == 5'h0 ? 5'h1 : _GEN_2; // @[BFS.scala 949:73 BFS.scala 950:12]
  wire [4:0] _GEN_4 = status == 5'h11 & tier_status_0 == 5'h0 ? 5'h2 : _GEN_3; // @[BFS.scala 947:73 BFS.scala 948:12]
  wire [4:0] _GEN_5 = io_signal & status == 5'h8 ? _GEN_1 : _GEN_4; // @[BFS.scala 941:55]
  wire [4:0] _GEN_6 = status == 5'h6 & io_cacheable_out_valid & io_cacheable_out_ready ? 5'h8 : _GEN_5; // @[BFS.scala 939:92 BFS.scala 940:12]
  wire [4:0] _GEN_7 = status == 5'h1 & tier_counter_1 == 32'h0 ? 5'h6 : _GEN_6; // @[BFS.scala 937:70 BFS.scala 938:12]
  wire [4:0] _GEN_8 = io_signal & status == 5'h7 ? _GEN_0 : _GEN_7; // @[BFS.scala 931:55]
  wire  next_tier_mask_hi = _T_2 | _T_5 | _T_8 | _T_23; // @[BFS.scala 955:115]
  wire  next_tier_mask_lo = _T_11 | _T_14 | _T_17 | _T_20; // @[BFS.scala 956:94]
  wire [1:0] next_tier_mask = {next_tier_mask_hi,next_tier_mask_lo}; // @[Cat.scala 30:58]
  reg [63:0] tier_base_addr_0; // @[BFS.scala 958:31]
  reg [63:0] tier_base_addr_1; // @[BFS.scala 958:31]
  wire  _step_fin_T_2 = _T_8 | _T_17; // @[BFS.scala 959:60]
  wire  step_fin = io_signal & (_T_8 | _T_17); // @[BFS.scala 959:28]
  wire  _axi_aw_valid_T_1 = tier_status_0 == 5'h3; // @[BFS.scala 1045:57]
  wire  _axi_aw_valid_T_2 = tier_status_1 == 5'h3; // @[BFS.scala 1045:90]
  wire  axi_aw_valid = next_tier_mask[0] ? tier_status_0 == 5'h3 : tier_status_1 == 5'h3; // @[BFS.scala 1045:22]
  wire [63:0] _tier_base_addr_0_T_1 = tier_base_addr_0 + 64'h400; // @[BFS.scala 965:16]
  wire  _T_35 = ~next_tier_mask[0]; // @[BFS.scala 966:18]
  wire  _axi_ar_valid_T_1 = tier_status_1 == 5'h4; // @[BFS.scala 1052:57]
  wire  _axi_ar_valid_T_2 = tier_status_0 == 5'h4; // @[BFS.scala 1052:89]
  wire  axi_ar_valid = next_tier_mask[0] ? tier_status_1 == 5'h4 : tier_status_0 == 5'h4; // @[BFS.scala 1052:22]
  wire [63:0] _tier_base_addr_1_T_1 = tier_base_addr_1 + 64'h400; // @[BFS.scala 965:16]
  wire  _T_49 = ~next_tier_mask[1]; // @[BFS.scala 966:18]
  wire  _T_55 = io_cacheable_in_0_ready & io_cacheable_in_0_valid; // @[BFS.scala 973:72]
  wire  _T_56 = io_cacheable_in_1_ready & io_cacheable_in_1_valid; // @[BFS.scala 973:72]
  wire  _T_57 = io_cacheable_in_2_ready & io_cacheable_in_2_valid; // @[BFS.scala 973:72]
  wire  _T_58 = io_cacheable_in_3_ready & io_cacheable_in_3_valid; // @[BFS.scala 973:72]
  wire  _T_59 = io_cacheable_in_4_ready & io_cacheable_in_4_valid; // @[BFS.scala 973:72]
  wire  _T_60 = io_cacheable_in_5_ready & io_cacheable_in_5_valid; // @[BFS.scala 973:72]
  wire  _T_61 = io_cacheable_in_6_ready & io_cacheable_in_6_valid; // @[BFS.scala 973:72]
  wire  _T_62 = io_cacheable_in_7_ready & io_cacheable_in_7_valid; // @[BFS.scala 973:72]
  wire  _T_63 = io_cacheable_in_8_ready & io_cacheable_in_8_valid; // @[BFS.scala 973:72]
  wire  _T_64 = io_cacheable_in_9_ready & io_cacheable_in_9_valid; // @[BFS.scala 973:72]
  wire  _T_65 = io_cacheable_in_10_ready & io_cacheable_in_10_valid; // @[BFS.scala 973:72]
  wire  _T_66 = io_cacheable_in_11_ready & io_cacheable_in_11_valid; // @[BFS.scala 973:72]
  wire  _T_67 = io_cacheable_in_12_ready & io_cacheable_in_12_valid; // @[BFS.scala 973:72]
  wire  _T_68 = io_cacheable_in_13_ready & io_cacheable_in_13_valid; // @[BFS.scala 973:72]
  wire  _T_69 = io_cacheable_in_14_ready & io_cacheable_in_14_valid; // @[BFS.scala 973:72]
  wire  _T_70 = io_cacheable_in_15_ready & io_cacheable_in_15_valid; // @[BFS.scala 973:72]
  wire  _T_85 = io_cacheable_in_0_ready & io_cacheable_in_0_valid | io_cacheable_in_1_ready & io_cacheable_in_1_valid |
    io_cacheable_in_2_ready & io_cacheable_in_2_valid | io_cacheable_in_3_ready & io_cacheable_in_3_valid |
    io_cacheable_in_4_ready & io_cacheable_in_4_valid | io_cacheable_in_5_ready & io_cacheable_in_5_valid |
    io_cacheable_in_6_ready & io_cacheable_in_6_valid | io_cacheable_in_7_ready & io_cacheable_in_7_valid |
    io_cacheable_in_8_ready & io_cacheable_in_8_valid | io_cacheable_in_9_ready & io_cacheable_in_9_valid |
    io_cacheable_in_10_ready & io_cacheable_in_10_valid | io_cacheable_in_11_ready & io_cacheable_in_11_valid |
    io_cacheable_in_12_ready & io_cacheable_in_12_valid | io_cacheable_in_13_ready & io_cacheable_in_13_valid |
    io_cacheable_in_14_ready & io_cacheable_in_14_valid | _T_70; // @[BFS.scala 973:93]
  wire [5:0] _tier_counter_0_WIRE = {{5'd0}, _T_55}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_WIRE_1 = {{5'd0}, _T_56}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_17 = _tier_counter_0_WIRE + _tier_counter_0_WIRE_1; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_2 = {{5'd0}, _T_57}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_19 = _tier_counter_0_T_17 + _tier_counter_0_WIRE_2; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_3 = {{5'd0}, _T_58}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_21 = _tier_counter_0_T_19 + _tier_counter_0_WIRE_3; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_4 = {{5'd0}, _T_59}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_23 = _tier_counter_0_T_21 + _tier_counter_0_WIRE_4; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_5 = {{5'd0}, _T_60}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_25 = _tier_counter_0_T_23 + _tier_counter_0_WIRE_5; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_6 = {{5'd0}, _T_61}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_27 = _tier_counter_0_T_25 + _tier_counter_0_WIRE_6; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_7 = {{5'd0}, _T_62}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_29 = _tier_counter_0_T_27 + _tier_counter_0_WIRE_7; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_8 = {{5'd0}, _T_63}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_31 = _tier_counter_0_T_29 + _tier_counter_0_WIRE_8; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_9 = {{5'd0}, _T_64}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_33 = _tier_counter_0_T_31 + _tier_counter_0_WIRE_9; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_10 = {{5'd0}, _T_65}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_35 = _tier_counter_0_T_33 + _tier_counter_0_WIRE_10; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_11 = {{5'd0}, _T_66}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_37 = _tier_counter_0_T_35 + _tier_counter_0_WIRE_11; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_12 = {{5'd0}, _T_67}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_39 = _tier_counter_0_T_37 + _tier_counter_0_WIRE_12; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_13 = {{5'd0}, _T_68}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_41 = _tier_counter_0_T_39 + _tier_counter_0_WIRE_13; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_14 = {{5'd0}, _T_69}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_43 = _tier_counter_0_T_41 + _tier_counter_0_WIRE_14; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_15 = {{5'd0}, _T_70}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_45 = _tier_counter_0_T_43 + _tier_counter_0_WIRE_15; // @[BFS.scala 974:100]
  wire [31:0] _GEN_36 = {{26'd0}, _tier_counter_0_T_45}; // @[BFS.scala 974:16]
  wire [31:0] _tier_counter_0_T_47 = tier_counter_0 + _GEN_36; // @[BFS.scala 974:16]
  wire [31:0] _tier_counter_0_T_50 = tier_counter_0 - 32'h10; // @[BFS.scala 976:59]
  wire [31:0] _GEN_37 = {{23'd0}, tier_fifo_0_io_out_data_count}; // @[BFS.scala 976:69]
  wire [31:0] _tier_counter_0_T_52 = tier_counter_0 - _GEN_37; // @[BFS.scala 976:69]
  wire [31:0] _tier_counter_1_T_47 = tier_counter_1 + _GEN_36; // @[BFS.scala 974:16]
  wire [31:0] _tier_counter_1_T_50 = tier_counter_1 - 32'h10; // @[BFS.scala 976:59]
  wire [31:0] _GEN_39 = {{23'd0}, tier_fifo_1_io_out_data_count}; // @[BFS.scala 976:69]
  wire [31:0] _tier_counter_1_T_52 = tier_counter_1 - _GEN_39; // @[BFS.scala 976:69]
  wire  _T_134 = tier_fifo_0_io_out_data_count == 9'h0; // @[BFS.scala 818:23]
  wire  _T_149 = tier_status_0 == 5'h9; // @[BFS.scala 1007:20]
  reg [7:0] wcount; // @[BFS.scala 1033:23]
  wire  axi_w_bits_wlast = wcount == 8'h1; // @[BFS.scala 1055:30]
  wire [4:0] _GEN_22 = tier_status_0 == 5'h9 & axi_w_bits_wlast & io_ddr_out_0_w_ready ? 5'h0 : tier_status_0; // @[BFS.scala 1007:94 BFS.scala 1008:11 BFS.scala 923:28]
  wire [4:0] _GEN_23 = tier_status_0 == 5'h10 & io_ddr_out_0_r_bits_rlast & io_ddr_out_0_r_valid ? 5'h0 : _GEN_22; // @[BFS.scala 1005:99 BFS.scala 1006:11]
  wire [4:0] _GEN_24 = _axi_ar_valid_T_2 & io_ddr_out_0_ar_ready ? 5'h10 : _GEN_23; // @[BFS.scala 1003:52 BFS.scala 1004:11]
  wire  _T_160 = tier_fifo_1_io_out_data_count == 9'h0; // @[BFS.scala 818:23]
  wire  _T_175 = tier_status_1 == 5'h9; // @[BFS.scala 1007:20]
  wire [4:0] _GEN_28 = tier_status_1 == 5'h9 & axi_w_bits_wlast & io_ddr_out_0_w_ready ? 5'h0 : tier_status_1; // @[BFS.scala 1007:94 BFS.scala 1008:11 BFS.scala 923:28]
  wire [4:0] _GEN_29 = tier_status_1 == 5'h10 & io_ddr_out_0_r_bits_rlast & io_ddr_out_0_r_valid ? 5'h0 : _GEN_28; // @[BFS.scala 1005:99 BFS.scala 1006:11]
  wire [4:0] _GEN_30 = _axi_ar_valid_T_1 & io_ddr_out_0_ar_ready ? 5'h10 : _GEN_29; // @[BFS.scala 1003:52 BFS.scala 1004:11]
  wire  _io_cacheable_out_valid_T_2 = tier_fifo_1_io_out_valid | _T_14; // @[BFS.scala 1020:57]
  wire  _io_cacheable_out_valid_T_5 = tier_fifo_0_io_out_valid | _T_5; // @[BFS.scala 1021:57]
  wire [511:0] _io_cacheable_out_bits_tdata_T_4 = next_tier_mask[1] ? tier_fifo_0_io_out_dout : 512'h0; // @[Mux.scala 98:16]
  wire [511:0] _io_cacheable_out_bits_tdata_T_5 = next_tier_mask[0] ? tier_fifo_1_io_out_dout :
    _io_cacheable_out_bits_tdata_T_4; // @[Mux.scala 98:16]
  wire [511:0] _io_cacheable_out_bits_tdata_T_6 = _T_14 ? 512'h80000000 : _io_cacheable_out_bits_tdata_T_5; // @[Mux.scala 98:16]
  wire  _io_cacheable_out_bits_tkeep_T_6 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h0 :
    tier_fifo_0_io_out_data_count > 9'h0; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_10 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h1 :
    tier_fifo_0_io_out_data_count > 9'h1; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_14 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h2 :
    tier_fifo_0_io_out_data_count > 9'h2; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_18 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h3 :
    tier_fifo_0_io_out_data_count > 9'h3; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_22 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h4 :
    tier_fifo_0_io_out_data_count > 9'h4; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_26 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h5 :
    tier_fifo_0_io_out_data_count > 9'h5; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_30 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h6 :
    tier_fifo_0_io_out_data_count > 9'h6; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_34 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h7 :
    tier_fifo_0_io_out_data_count > 9'h7; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_38 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h8 :
    tier_fifo_0_io_out_data_count > 9'h8; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_42 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h9 :
    tier_fifo_0_io_out_data_count > 9'h9; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_46 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'ha :
    tier_fifo_0_io_out_data_count > 9'ha; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_50 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'hb :
    tier_fifo_0_io_out_data_count > 9'hb; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_54 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'hc :
    tier_fifo_0_io_out_data_count > 9'hc; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_58 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'hd :
    tier_fifo_0_io_out_data_count > 9'hd; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_62 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'he :
    tier_fifo_0_io_out_data_count > 9'he; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_66 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'hf :
    tier_fifo_0_io_out_data_count > 9'hf; // @[BFS.scala 1029:15]
  wire [7:0] io_cacheable_out_bits_tkeep_lo = {_io_cacheable_out_bits_tkeep_T_34,_io_cacheable_out_bits_tkeep_T_30,
    _io_cacheable_out_bits_tkeep_T_26,_io_cacheable_out_bits_tkeep_T_22,_io_cacheable_out_bits_tkeep_T_18,
    _io_cacheable_out_bits_tkeep_T_14,_io_cacheable_out_bits_tkeep_T_10,_io_cacheable_out_bits_tkeep_T_6}; // @[BFS.scala 1030:14]
  wire [15:0] _io_cacheable_out_bits_tkeep_T_67 = {_io_cacheable_out_bits_tkeep_T_66,_io_cacheable_out_bits_tkeep_T_62,
    _io_cacheable_out_bits_tkeep_T_58,_io_cacheable_out_bits_tkeep_T_54,_io_cacheable_out_bits_tkeep_T_50,
    _io_cacheable_out_bits_tkeep_T_46,_io_cacheable_out_bits_tkeep_T_42,_io_cacheable_out_bits_tkeep_T_38,
    io_cacheable_out_bits_tkeep_lo}; // @[BFS.scala 1030:14]
  wire  axi_w_valid = next_tier_mask[0] ? _T_149 : _T_175; // @[BFS.scala 1054:21]
  wire [7:0] _wcount_T_1 = wcount - 8'h1; // @[BFS.scala 1037:22]
  multi_channel_fifo tier_fifo_0 ( // @[BFS.scala 903:46]
    .clock(tier_fifo_0_clock),
    .reset(tier_fifo_0_reset),
    .io_in_0_ready(tier_fifo_0_io_in_0_ready),
    .io_in_0_valid(tier_fifo_0_io_in_0_valid),
    .io_in_0_bits_tdata(tier_fifo_0_io_in_0_bits_tdata),
    .io_in_1_ready(tier_fifo_0_io_in_1_ready),
    .io_in_1_valid(tier_fifo_0_io_in_1_valid),
    .io_in_1_bits_tdata(tier_fifo_0_io_in_1_bits_tdata),
    .io_in_2_ready(tier_fifo_0_io_in_2_ready),
    .io_in_2_valid(tier_fifo_0_io_in_2_valid),
    .io_in_2_bits_tdata(tier_fifo_0_io_in_2_bits_tdata),
    .io_in_3_ready(tier_fifo_0_io_in_3_ready),
    .io_in_3_valid(tier_fifo_0_io_in_3_valid),
    .io_in_3_bits_tdata(tier_fifo_0_io_in_3_bits_tdata),
    .io_in_4_ready(tier_fifo_0_io_in_4_ready),
    .io_in_4_valid(tier_fifo_0_io_in_4_valid),
    .io_in_4_bits_tdata(tier_fifo_0_io_in_4_bits_tdata),
    .io_in_5_ready(tier_fifo_0_io_in_5_ready),
    .io_in_5_valid(tier_fifo_0_io_in_5_valid),
    .io_in_5_bits_tdata(tier_fifo_0_io_in_5_bits_tdata),
    .io_in_6_ready(tier_fifo_0_io_in_6_ready),
    .io_in_6_valid(tier_fifo_0_io_in_6_valid),
    .io_in_6_bits_tdata(tier_fifo_0_io_in_6_bits_tdata),
    .io_in_7_ready(tier_fifo_0_io_in_7_ready),
    .io_in_7_valid(tier_fifo_0_io_in_7_valid),
    .io_in_7_bits_tdata(tier_fifo_0_io_in_7_bits_tdata),
    .io_in_8_ready(tier_fifo_0_io_in_8_ready),
    .io_in_8_valid(tier_fifo_0_io_in_8_valid),
    .io_in_8_bits_tdata(tier_fifo_0_io_in_8_bits_tdata),
    .io_in_9_ready(tier_fifo_0_io_in_9_ready),
    .io_in_9_valid(tier_fifo_0_io_in_9_valid),
    .io_in_9_bits_tdata(tier_fifo_0_io_in_9_bits_tdata),
    .io_in_10_ready(tier_fifo_0_io_in_10_ready),
    .io_in_10_valid(tier_fifo_0_io_in_10_valid),
    .io_in_10_bits_tdata(tier_fifo_0_io_in_10_bits_tdata),
    .io_in_11_ready(tier_fifo_0_io_in_11_ready),
    .io_in_11_valid(tier_fifo_0_io_in_11_valid),
    .io_in_11_bits_tdata(tier_fifo_0_io_in_11_bits_tdata),
    .io_in_12_ready(tier_fifo_0_io_in_12_ready),
    .io_in_12_valid(tier_fifo_0_io_in_12_valid),
    .io_in_12_bits_tdata(tier_fifo_0_io_in_12_bits_tdata),
    .io_in_13_ready(tier_fifo_0_io_in_13_ready),
    .io_in_13_valid(tier_fifo_0_io_in_13_valid),
    .io_in_13_bits_tdata(tier_fifo_0_io_in_13_bits_tdata),
    .io_in_14_ready(tier_fifo_0_io_in_14_ready),
    .io_in_14_valid(tier_fifo_0_io_in_14_valid),
    .io_in_14_bits_tdata(tier_fifo_0_io_in_14_bits_tdata),
    .io_in_15_ready(tier_fifo_0_io_in_15_ready),
    .io_in_15_valid(tier_fifo_0_io_in_15_valid),
    .io_in_15_bits_tdata(tier_fifo_0_io_in_15_bits_tdata),
    .io_out_full(tier_fifo_0_io_out_full),
    .io_out_din(tier_fifo_0_io_out_din),
    .io_out_wr_en(tier_fifo_0_io_out_wr_en),
    .io_out_dout(tier_fifo_0_io_out_dout),
    .io_out_rd_en(tier_fifo_0_io_out_rd_en),
    .io_out_data_count(tier_fifo_0_io_out_data_count),
    .io_out_valid(tier_fifo_0_io_out_valid),
    .io_flush(tier_fifo_0_io_flush),
    .io_is_current_tier(tier_fifo_0_io_is_current_tier)
  );
  multi_channel_fifo tier_fifo_1 ( // @[BFS.scala 903:46]
    .clock(tier_fifo_1_clock),
    .reset(tier_fifo_1_reset),
    .io_in_0_ready(tier_fifo_1_io_in_0_ready),
    .io_in_0_valid(tier_fifo_1_io_in_0_valid),
    .io_in_0_bits_tdata(tier_fifo_1_io_in_0_bits_tdata),
    .io_in_1_ready(tier_fifo_1_io_in_1_ready),
    .io_in_1_valid(tier_fifo_1_io_in_1_valid),
    .io_in_1_bits_tdata(tier_fifo_1_io_in_1_bits_tdata),
    .io_in_2_ready(tier_fifo_1_io_in_2_ready),
    .io_in_2_valid(tier_fifo_1_io_in_2_valid),
    .io_in_2_bits_tdata(tier_fifo_1_io_in_2_bits_tdata),
    .io_in_3_ready(tier_fifo_1_io_in_3_ready),
    .io_in_3_valid(tier_fifo_1_io_in_3_valid),
    .io_in_3_bits_tdata(tier_fifo_1_io_in_3_bits_tdata),
    .io_in_4_ready(tier_fifo_1_io_in_4_ready),
    .io_in_4_valid(tier_fifo_1_io_in_4_valid),
    .io_in_4_bits_tdata(tier_fifo_1_io_in_4_bits_tdata),
    .io_in_5_ready(tier_fifo_1_io_in_5_ready),
    .io_in_5_valid(tier_fifo_1_io_in_5_valid),
    .io_in_5_bits_tdata(tier_fifo_1_io_in_5_bits_tdata),
    .io_in_6_ready(tier_fifo_1_io_in_6_ready),
    .io_in_6_valid(tier_fifo_1_io_in_6_valid),
    .io_in_6_bits_tdata(tier_fifo_1_io_in_6_bits_tdata),
    .io_in_7_ready(tier_fifo_1_io_in_7_ready),
    .io_in_7_valid(tier_fifo_1_io_in_7_valid),
    .io_in_7_bits_tdata(tier_fifo_1_io_in_7_bits_tdata),
    .io_in_8_ready(tier_fifo_1_io_in_8_ready),
    .io_in_8_valid(tier_fifo_1_io_in_8_valid),
    .io_in_8_bits_tdata(tier_fifo_1_io_in_8_bits_tdata),
    .io_in_9_ready(tier_fifo_1_io_in_9_ready),
    .io_in_9_valid(tier_fifo_1_io_in_9_valid),
    .io_in_9_bits_tdata(tier_fifo_1_io_in_9_bits_tdata),
    .io_in_10_ready(tier_fifo_1_io_in_10_ready),
    .io_in_10_valid(tier_fifo_1_io_in_10_valid),
    .io_in_10_bits_tdata(tier_fifo_1_io_in_10_bits_tdata),
    .io_in_11_ready(tier_fifo_1_io_in_11_ready),
    .io_in_11_valid(tier_fifo_1_io_in_11_valid),
    .io_in_11_bits_tdata(tier_fifo_1_io_in_11_bits_tdata),
    .io_in_12_ready(tier_fifo_1_io_in_12_ready),
    .io_in_12_valid(tier_fifo_1_io_in_12_valid),
    .io_in_12_bits_tdata(tier_fifo_1_io_in_12_bits_tdata),
    .io_in_13_ready(tier_fifo_1_io_in_13_ready),
    .io_in_13_valid(tier_fifo_1_io_in_13_valid),
    .io_in_13_bits_tdata(tier_fifo_1_io_in_13_bits_tdata),
    .io_in_14_ready(tier_fifo_1_io_in_14_ready),
    .io_in_14_valid(tier_fifo_1_io_in_14_valid),
    .io_in_14_bits_tdata(tier_fifo_1_io_in_14_bits_tdata),
    .io_in_15_ready(tier_fifo_1_io_in_15_ready),
    .io_in_15_valid(tier_fifo_1_io_in_15_valid),
    .io_in_15_bits_tdata(tier_fifo_1_io_in_15_bits_tdata),
    .io_out_full(tier_fifo_1_io_out_full),
    .io_out_din(tier_fifo_1_io_out_din),
    .io_out_wr_en(tier_fifo_1_io_out_wr_en),
    .io_out_dout(tier_fifo_1_io_out_dout),
    .io_out_rd_en(tier_fifo_1_io_out_rd_en),
    .io_out_data_count(tier_fifo_1_io_out_data_count),
    .io_out_valid(tier_fifo_1_io_out_valid),
    .io_flush(tier_fifo_1_io_flush),
    .io_is_current_tier(tier_fifo_1_io_is_current_tier)
  );
  assign io_cacheable_out_valid = next_tier_mask[0] ? _io_cacheable_out_valid_T_2 : next_tier_mask[1] &
    _io_cacheable_out_valid_T_5; // @[Mux.scala 98:16]
  assign io_cacheable_out_bits_tdata = _T_5 ? 512'h80000000 : _io_cacheable_out_bits_tdata_T_6; // @[Mux.scala 98:16]
  assign io_cacheable_out_bits_tkeep = _T_5 | _T_14 ? 16'h1 : _io_cacheable_out_bits_tkeep_T_67; // @[BFS.scala 1027:37]
  assign io_cacheable_in_0_ready = next_tier_mask[0] ? tier_fifo_0_io_in_0_ready : tier_fifo_1_io_in_0_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_1_ready = next_tier_mask[0] ? tier_fifo_0_io_in_1_ready : tier_fifo_1_io_in_1_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_2_ready = next_tier_mask[0] ? tier_fifo_0_io_in_2_ready : tier_fifo_1_io_in_2_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_3_ready = next_tier_mask[0] ? tier_fifo_0_io_in_3_ready : tier_fifo_1_io_in_3_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_4_ready = next_tier_mask[0] ? tier_fifo_0_io_in_4_ready : tier_fifo_1_io_in_4_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_5_ready = next_tier_mask[0] ? tier_fifo_0_io_in_5_ready : tier_fifo_1_io_in_5_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_6_ready = next_tier_mask[0] ? tier_fifo_0_io_in_6_ready : tier_fifo_1_io_in_6_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_7_ready = next_tier_mask[0] ? tier_fifo_0_io_in_7_ready : tier_fifo_1_io_in_7_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_8_ready = next_tier_mask[0] ? tier_fifo_0_io_in_8_ready : tier_fifo_1_io_in_8_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_9_ready = next_tier_mask[0] ? tier_fifo_0_io_in_9_ready : tier_fifo_1_io_in_9_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_10_ready = next_tier_mask[0] ? tier_fifo_0_io_in_10_ready : tier_fifo_1_io_in_10_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_11_ready = next_tier_mask[0] ? tier_fifo_0_io_in_11_ready : tier_fifo_1_io_in_11_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_12_ready = next_tier_mask[0] ? tier_fifo_0_io_in_12_ready : tier_fifo_1_io_in_12_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_13_ready = next_tier_mask[0] ? tier_fifo_0_io_in_13_ready : tier_fifo_1_io_in_13_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_14_ready = next_tier_mask[0] ? tier_fifo_0_io_in_14_ready : tier_fifo_1_io_in_14_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_15_ready = next_tier_mask[0] ? tier_fifo_0_io_in_15_ready : tier_fifo_1_io_in_15_ready; // @[BFS.scala 1015:22]
  assign io_non_cacheable_in_aw_ready = io_ddr_out_1_aw_ready; // @[BFS.scala 1061:17]
  assign io_non_cacheable_in_w_ready = io_ddr_out_1_w_ready; // @[BFS.scala 1061:17]
  assign io_ddr_out_0_aw_valid = next_tier_mask[0] ? tier_status_0 == 5'h3 : tier_status_1 == 5'h3; // @[BFS.scala 1045:22]
  assign io_ddr_out_0_aw_bits_awaddr = next_tier_mask[0] ? tier_base_addr_0 : tier_base_addr_1; // @[BFS.scala 1039:28]
  assign io_ddr_out_0_ar_valid = next_tier_mask[0] ? tier_status_1 == 5'h4 : tier_status_0 == 5'h4; // @[BFS.scala 1052:22]
  assign io_ddr_out_0_ar_bits_araddr = next_tier_mask[0] ? tier_base_addr_1 : tier_base_addr_0; // @[BFS.scala 1046:28]
  assign io_ddr_out_0_w_valid = next_tier_mask[0] ? _T_149 : _T_175; // @[BFS.scala 1054:21]
  assign io_ddr_out_0_w_bits_wdata = next_tier_mask[0] ? tier_fifo_0_io_out_dout : tier_fifo_1_io_out_dout; // @[BFS.scala 1053:26]
  assign io_ddr_out_0_w_bits_wlast = wcount == 8'h1; // @[BFS.scala 1055:30]
  assign io_ddr_out_1_aw_valid = io_non_cacheable_in_aw_valid; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_aw_bits_awaddr = io_non_cacheable_in_aw_bits_awaddr; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_aw_bits_awid = io_non_cacheable_in_aw_bits_awid; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_w_valid = io_non_cacheable_in_w_valid; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_w_bits_wdata = io_non_cacheable_in_w_bits_wdata; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_w_bits_wstrb = io_non_cacheable_in_w_bits_wstrb; // @[BFS.scala 1061:17]
  assign io_unvisited_size = next_tier_mask[0] ? tier_counter_0 : tier_counter_1; // @[BFS.scala 1018:27]
  assign tier_fifo_0_clock = clock;
  assign tier_fifo_0_reset = reset;
  assign tier_fifo_0_io_in_0_valid = next_tier_mask[0] & io_cacheable_in_0_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_0_bits_tdata = next_tier_mask[0] ? io_cacheable_in_0_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_1_valid = next_tier_mask[0] & io_cacheable_in_1_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_1_bits_tdata = next_tier_mask[0] ? io_cacheable_in_1_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_2_valid = next_tier_mask[0] & io_cacheable_in_2_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_2_bits_tdata = next_tier_mask[0] ? io_cacheable_in_2_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_3_valid = next_tier_mask[0] & io_cacheable_in_3_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_3_bits_tdata = next_tier_mask[0] ? io_cacheable_in_3_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_4_valid = next_tier_mask[0] & io_cacheable_in_4_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_4_bits_tdata = next_tier_mask[0] ? io_cacheable_in_4_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_5_valid = next_tier_mask[0] & io_cacheable_in_5_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_5_bits_tdata = next_tier_mask[0] ? io_cacheable_in_5_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_6_valid = next_tier_mask[0] & io_cacheable_in_6_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_6_bits_tdata = next_tier_mask[0] ? io_cacheable_in_6_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_7_valid = next_tier_mask[0] & io_cacheable_in_7_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_7_bits_tdata = next_tier_mask[0] ? io_cacheable_in_7_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_8_valid = next_tier_mask[0] & io_cacheable_in_8_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_8_bits_tdata = next_tier_mask[0] ? io_cacheable_in_8_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_9_valid = next_tier_mask[0] & io_cacheable_in_9_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_9_bits_tdata = next_tier_mask[0] ? io_cacheable_in_9_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_10_valid = next_tier_mask[0] & io_cacheable_in_10_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_10_bits_tdata = next_tier_mask[0] ? io_cacheable_in_10_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_11_valid = next_tier_mask[0] & io_cacheable_in_11_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_11_bits_tdata = next_tier_mask[0] ? io_cacheable_in_11_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_12_valid = next_tier_mask[0] & io_cacheable_in_12_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_12_bits_tdata = next_tier_mask[0] ? io_cacheable_in_12_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_13_valid = next_tier_mask[0] & io_cacheable_in_13_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_13_bits_tdata = next_tier_mask[0] ? io_cacheable_in_13_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_14_valid = next_tier_mask[0] & io_cacheable_in_14_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_14_bits_tdata = next_tier_mask[0] ? io_cacheable_in_14_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_15_valid = next_tier_mask[0] & io_cacheable_in_15_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_15_bits_tdata = next_tier_mask[0] ? io_cacheable_in_15_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_out_din = next_tier_mask[0] ? 512'h0 : io_ddr_out_0_r_bits_rdata; // @[BFS.scala 984:26]
  assign tier_fifo_0_io_out_wr_en = next_tier_mask[0] ? 1'h0 : io_ddr_out_0_r_valid; // @[BFS.scala 983:28]
  assign tier_fifo_0_io_out_rd_en = next_tier_mask[0] ? io_ddr_out_0_w_ready : io_cacheable_out_ready; // @[BFS.scala 982:28]
  assign tier_fifo_0_io_flush = io_signal & _step_fin_T_2; // @[BFS.scala 985:31]
  assign tier_fifo_0_io_is_current_tier = ~next_tier_mask[0]; // @[BFS.scala 992:31]
  assign tier_fifo_1_clock = clock;
  assign tier_fifo_1_reset = reset;
  assign tier_fifo_1_io_in_0_valid = next_tier_mask[1] & io_cacheable_in_0_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_0_bits_tdata = next_tier_mask[1] ? io_cacheable_in_0_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_1_valid = next_tier_mask[1] & io_cacheable_in_1_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_1_bits_tdata = next_tier_mask[1] ? io_cacheable_in_1_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_2_valid = next_tier_mask[1] & io_cacheable_in_2_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_2_bits_tdata = next_tier_mask[1] ? io_cacheable_in_2_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_3_valid = next_tier_mask[1] & io_cacheable_in_3_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_3_bits_tdata = next_tier_mask[1] ? io_cacheable_in_3_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_4_valid = next_tier_mask[1] & io_cacheable_in_4_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_4_bits_tdata = next_tier_mask[1] ? io_cacheable_in_4_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_5_valid = next_tier_mask[1] & io_cacheable_in_5_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_5_bits_tdata = next_tier_mask[1] ? io_cacheable_in_5_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_6_valid = next_tier_mask[1] & io_cacheable_in_6_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_6_bits_tdata = next_tier_mask[1] ? io_cacheable_in_6_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_7_valid = next_tier_mask[1] & io_cacheable_in_7_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_7_bits_tdata = next_tier_mask[1] ? io_cacheable_in_7_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_8_valid = next_tier_mask[1] & io_cacheable_in_8_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_8_bits_tdata = next_tier_mask[1] ? io_cacheable_in_8_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_9_valid = next_tier_mask[1] & io_cacheable_in_9_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_9_bits_tdata = next_tier_mask[1] ? io_cacheable_in_9_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_10_valid = next_tier_mask[1] & io_cacheable_in_10_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_10_bits_tdata = next_tier_mask[1] ? io_cacheable_in_10_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_11_valid = next_tier_mask[1] & io_cacheable_in_11_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_11_bits_tdata = next_tier_mask[1] ? io_cacheable_in_11_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_12_valid = next_tier_mask[1] & io_cacheable_in_12_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_12_bits_tdata = next_tier_mask[1] ? io_cacheable_in_12_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_13_valid = next_tier_mask[1] & io_cacheable_in_13_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_13_bits_tdata = next_tier_mask[1] ? io_cacheable_in_13_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_14_valid = next_tier_mask[1] & io_cacheable_in_14_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_14_bits_tdata = next_tier_mask[1] ? io_cacheable_in_14_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_15_valid = next_tier_mask[1] & io_cacheable_in_15_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_15_bits_tdata = next_tier_mask[1] ? io_cacheable_in_15_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_out_din = next_tier_mask[1] ? 512'h0 : io_ddr_out_0_r_bits_rdata; // @[BFS.scala 984:26]
  assign tier_fifo_1_io_out_wr_en = next_tier_mask[1] ? 1'h0 : io_ddr_out_0_r_valid; // @[BFS.scala 983:28]
  assign tier_fifo_1_io_out_rd_en = next_tier_mask[1] ? io_ddr_out_0_w_ready : io_cacheable_out_ready; // @[BFS.scala 982:28]
  assign tier_fifo_1_io_flush = io_signal & _step_fin_T_2; // @[BFS.scala 985:31]
  assign tier_fifo_1_io_is_current_tier = ~next_tier_mask[1]; // @[BFS.scala 992:31]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 904:29]
      tier_counter_0 <= 32'h0; // @[BFS.scala 904:29]
    end else if (next_tier_mask[0] & _T_85) begin // @[BFS.scala 973:97]
      tier_counter_0 <= _tier_counter_0_T_47; // @[BFS.scala 974:11]
    end else if (_T_35 & io_cacheable_out_ready & io_cacheable_out_valid) begin // @[BFS.scala 975:89]
      if (tier_fifo_0_io_out_data_count > 9'h10) begin // @[BFS.scala 976:17]
        tier_counter_0 <= _tier_counter_0_T_50;
      end else begin
        tier_counter_0 <= _tier_counter_0_T_52;
      end
    end
    if (reset) begin // @[BFS.scala 904:29]
      tier_counter_1 <= 32'h0; // @[BFS.scala 904:29]
    end else if (next_tier_mask[1] & _T_85) begin // @[BFS.scala 973:97]
      tier_counter_1 <= _tier_counter_1_T_47; // @[BFS.scala 974:11]
    end else if (_T_49 & io_cacheable_out_ready & io_cacheable_out_valid) begin // @[BFS.scala 975:89]
      if (tier_fifo_1_io_out_data_count > 9'h10) begin // @[BFS.scala 976:17]
        tier_counter_1 <= _tier_counter_1_T_50;
      end else begin
        tier_counter_1 <= _tier_counter_1_T_52;
      end
    end
    if (reset) begin // @[BFS.scala 922:23]
      status <= 5'h0; // @[BFS.scala 922:23]
    end else if (io_start & status == 5'h0) begin // @[BFS.scala 925:40]
      status <= 5'h2; // @[BFS.scala 926:12]
    end else if (status == 5'h2 & tier_counter_0 == 32'h0) begin // @[BFS.scala 927:70]
      status <= 5'h5; // @[BFS.scala 928:12]
    end else if (status == 5'h5 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 929:92]
      status <= 5'h7; // @[BFS.scala 930:12]
    end else begin
      status <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 923:28]
      tier_status_0 <= 5'h0; // @[BFS.scala 923:28]
    end else if (next_tier_mask[0] & tier_fifo_0_io_out_full & _T_21) begin // @[BFS.scala 997:76]
      tier_status_0 <= 5'h3; // @[BFS.scala 998:11]
    end else if (_T_35 & _T_134 & tier_counter_0 != 32'h0 & _T_21) begin // @[BFS.scala 999:109]
      tier_status_0 <= 5'h4; // @[BFS.scala 1000:11]
    end else if (_axi_aw_valid_T_1 & io_ddr_out_0_aw_ready) begin // @[BFS.scala 1001:53]
      tier_status_0 <= 5'h9; // @[BFS.scala 1002:11]
    end else begin
      tier_status_0 <= _GEN_24;
    end
    if (reset) begin // @[BFS.scala 923:28]
      tier_status_1 <= 5'h0; // @[BFS.scala 923:28]
    end else if (next_tier_mask[1] & tier_fifo_1_io_out_full & _T_24) begin // @[BFS.scala 997:76]
      tier_status_1 <= 5'h3; // @[BFS.scala 998:11]
    end else if (_T_49 & _T_160 & tier_counter_1 != 32'h0 & _T_24) begin // @[BFS.scala 999:109]
      tier_status_1 <= 5'h4; // @[BFS.scala 1000:11]
    end else if (_axi_aw_valid_T_2 & io_ddr_out_0_aw_ready) begin // @[BFS.scala 1001:53]
      tier_status_1 <= 5'h9; // @[BFS.scala 1002:11]
    end else begin
      tier_status_1 <= _GEN_30;
    end
    if (reset) begin // @[BFS.scala 958:31]
      tier_base_addr_0 <= 64'h0; // @[BFS.scala 958:31]
    end else if (_T_1 | step_fin) begin // @[BFS.scala 962:57]
      tier_base_addr_0 <= io_tiers_base_addr_0; // @[BFS.scala 963:11]
    end else if (next_tier_mask[0] & io_ddr_out_0_aw_ready & axi_aw_valid) begin // @[BFS.scala 964:86]
      tier_base_addr_0 <= _tier_base_addr_0_T_1; // @[BFS.scala 965:11]
    end else if (~next_tier_mask[0] & io_ddr_out_0_ar_ready & axi_ar_valid) begin // @[BFS.scala 966:87]
      tier_base_addr_0 <= _tier_base_addr_0_T_1; // @[BFS.scala 967:11]
    end
    if (reset) begin // @[BFS.scala 958:31]
      tier_base_addr_1 <= 64'h0; // @[BFS.scala 958:31]
    end else if (_T_1 | step_fin) begin // @[BFS.scala 962:57]
      tier_base_addr_1 <= io_tiers_base_addr_1; // @[BFS.scala 963:11]
    end else if (next_tier_mask[1] & io_ddr_out_0_aw_ready & axi_aw_valid) begin // @[BFS.scala 964:86]
      tier_base_addr_1 <= _tier_base_addr_1_T_1; // @[BFS.scala 965:11]
    end else if (~next_tier_mask[1] & io_ddr_out_0_ar_ready & axi_ar_valid) begin // @[BFS.scala 966:87]
      tier_base_addr_1 <= _tier_base_addr_1_T_1; // @[BFS.scala 967:11]
    end
    if (reset) begin // @[BFS.scala 1033:23]
      wcount <= 8'h0; // @[BFS.scala 1033:23]
    end else if (axi_aw_valid & io_ddr_out_0_aw_ready) begin // @[BFS.scala 1034:55]
      wcount <= 8'h10; // @[BFS.scala 1035:12]
    end else if (axi_w_valid & io_ddr_out_0_w_ready) begin // @[BFS.scala 1036:59]
      wcount <= _wcount_T_1; // @[BFS.scala 1037:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tier_counter_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  tier_counter_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  status = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  tier_status_0 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  tier_status_1 = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  tier_base_addr_0 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  tier_base_addr_1 = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  wcount = _RAND_7[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_arbitrator(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] data; // @[BFS.scala 237:21]
  reg [15:0] keep; // @[BFS.scala 238:21]
  wire  _T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 240:25]
  wire  _select_T_1 = |keep[0]; // @[BFS.scala 246:125]
  wire  _select_T_4 = |keep[1]; // @[BFS.scala 246:125]
  wire  _select_T_7 = |keep[2]; // @[BFS.scala 246:125]
  wire  _select_T_10 = |keep[3]; // @[BFS.scala 246:125]
  wire  _select_T_13 = |keep[4]; // @[BFS.scala 246:125]
  wire  _select_T_16 = |keep[5]; // @[BFS.scala 246:125]
  wire  _select_T_19 = |keep[6]; // @[BFS.scala 246:125]
  wire  _select_T_22 = |keep[7]; // @[BFS.scala 246:125]
  wire  _select_T_25 = |keep[8]; // @[BFS.scala 246:125]
  wire  _select_T_28 = |keep[9]; // @[BFS.scala 246:125]
  wire  _select_T_31 = |keep[10]; // @[BFS.scala 246:125]
  wire  _select_T_34 = |keep[11]; // @[BFS.scala 246:125]
  wire  _select_T_37 = |keep[12]; // @[BFS.scala 246:125]
  wire  _select_T_40 = |keep[13]; // @[BFS.scala 246:125]
  wire  _select_T_43 = |keep[14]; // @[BFS.scala 246:125]
  wire  _select_T_46 = |keep[15]; // @[BFS.scala 246:125]
  wire [30:0] _select_T_48 = _select_T_46 ? 31'h8000 : 31'h0; // @[Mux.scala 98:16]
  wire [30:0] _select_T_49 = _select_T_43 ? 31'h4000 : _select_T_48; // @[Mux.scala 98:16]
  wire [30:0] _select_T_50 = _select_T_40 ? 31'h2000 : _select_T_49; // @[Mux.scala 98:16]
  wire [30:0] _select_T_51 = _select_T_37 ? 31'h1000 : _select_T_50; // @[Mux.scala 98:16]
  wire [30:0] _select_T_52 = _select_T_34 ? 31'h800 : _select_T_51; // @[Mux.scala 98:16]
  wire [30:0] _select_T_53 = _select_T_31 ? 31'h400 : _select_T_52; // @[Mux.scala 98:16]
  wire [30:0] _select_T_54 = _select_T_28 ? 31'h200 : _select_T_53; // @[Mux.scala 98:16]
  wire [30:0] _select_T_55 = _select_T_25 ? 31'h100 : _select_T_54; // @[Mux.scala 98:16]
  wire [30:0] _select_T_56 = _select_T_22 ? 31'h80 : _select_T_55; // @[Mux.scala 98:16]
  wire [30:0] _select_T_57 = _select_T_19 ? 31'h40 : _select_T_56; // @[Mux.scala 98:16]
  wire [30:0] _select_T_58 = _select_T_16 ? 31'h20 : _select_T_57; // @[Mux.scala 98:16]
  wire [30:0] _select_T_59 = _select_T_13 ? 31'h10 : _select_T_58; // @[Mux.scala 98:16]
  wire [30:0] _select_T_60 = _select_T_10 ? 31'h8 : _select_T_59; // @[Mux.scala 98:16]
  wire [30:0] _select_T_61 = _select_T_7 ? 31'h4 : _select_T_60; // @[Mux.scala 98:16]
  wire [30:0] _select_T_62 = _select_T_4 ? 31'h2 : _select_T_61; // @[Mux.scala 98:16]
  wire [30:0] select = _select_T_1 ? 31'h1 : _select_T_62; // @[Mux.scala 98:16]
  wire [31:0] _io_ddr_out_bits_tdata_T_32 = select[0] ? data[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_33 = select[1] ? data[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_34 = select[2] ? data[95:64] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_35 = select[3] ? data[127:96] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_36 = select[4] ? data[159:128] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_37 = select[5] ? data[191:160] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_38 = select[6] ? data[223:192] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_39 = select[7] ? data[255:224] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_40 = select[8] ? data[287:256] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_41 = select[9] ? data[319:288] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_42 = select[10] ? data[351:320] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_43 = select[11] ? data[383:352] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_44 = select[12] ? data[415:384] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_45 = select[13] ? data[447:416] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_46 = select[14] ? data[479:448] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_47 = select[15] ? data[511:480] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_48 = _io_ddr_out_bits_tdata_T_32 | _io_ddr_out_bits_tdata_T_33; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_49 = _io_ddr_out_bits_tdata_T_48 | _io_ddr_out_bits_tdata_T_34; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_50 = _io_ddr_out_bits_tdata_T_49 | _io_ddr_out_bits_tdata_T_35; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_51 = _io_ddr_out_bits_tdata_T_50 | _io_ddr_out_bits_tdata_T_36; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_52 = _io_ddr_out_bits_tdata_T_51 | _io_ddr_out_bits_tdata_T_37; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_53 = _io_ddr_out_bits_tdata_T_52 | _io_ddr_out_bits_tdata_T_38; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_54 = _io_ddr_out_bits_tdata_T_53 | _io_ddr_out_bits_tdata_T_39; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_55 = _io_ddr_out_bits_tdata_T_54 | _io_ddr_out_bits_tdata_T_40; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_56 = _io_ddr_out_bits_tdata_T_55 | _io_ddr_out_bits_tdata_T_41; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_57 = _io_ddr_out_bits_tdata_T_56 | _io_ddr_out_bits_tdata_T_42; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_58 = _io_ddr_out_bits_tdata_T_57 | _io_ddr_out_bits_tdata_T_43; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_59 = _io_ddr_out_bits_tdata_T_58 | _io_ddr_out_bits_tdata_T_44; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_60 = _io_ddr_out_bits_tdata_T_59 | _io_ddr_out_bits_tdata_T_45; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_61 = _io_ddr_out_bits_tdata_T_60 | _io_ddr_out_bits_tdata_T_46; // @[Mux.scala 27:72]
  wire  next_keep_0 = select[0] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_1 = select[1] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_2 = select[2] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_3 = select[3] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_4 = select[4] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_5 = select[5] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_6 = select[6] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_7 = select[7] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_8 = select[8] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_9 = select[9] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_10 = select[10] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_11 = select[11] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_12 = select[12] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_13 = select[13] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_14 = select[14] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_15 = select[15] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire [7:0] keep_lo = {next_keep_7,next_keep_6,next_keep_5,next_keep_4,next_keep_3,next_keep_2,next_keep_1,next_keep_0}
    ; // @[BFS.scala 262:36]
  wire [15:0] _keep_T = {next_keep_15,next_keep_14,next_keep_13,next_keep_12,next_keep_11,next_keep_10,next_keep_9,
    next_keep_8,keep_lo}; // @[BFS.scala 262:36]
  wire [15:0] _keep_T_1 = keep & _keep_T; // @[BFS.scala 262:18]
  assign io_xbar_in_ready = ~(|keep); // @[BFS.scala 243:23]
  assign io_ddr_out_valid = |select; // @[BFS.scala 247:33]
  assign io_ddr_out_bits_tdata = _io_ddr_out_bits_tdata_T_61 | _io_ddr_out_bits_tdata_T_47; // @[Mux.scala 27:72]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 237:21]
      data <= 512'h0; // @[BFS.scala 237:21]
    end else if (io_xbar_in_valid & io_xbar_in_ready) begin // @[BFS.scala 240:45]
      data <= io_xbar_in_bits_tdata; // @[BFS.scala 241:10]
    end
    if (reset) begin // @[BFS.scala 238:21]
      keep <= 16'h0; // @[BFS.scala 238:21]
    end else if (_T) begin // @[BFS.scala 259:45]
      keep <= io_xbar_in_bits_tkeep; // @[BFS.scala 260:10]
    end else if (io_ddr_out_valid & io_ddr_out_ready) begin // @[BFS.scala 261:52]
      keep <= _keep_T_1; // @[BFS.scala 262:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  data = _RAND_0[511:0];
  _RAND_1 = {1{`RANDOM}};
  keep = _RAND_1[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pipeline_32(
  input         clock,
  input         reset,
  input         io_dout_ready,
  output        io_dout_valid,
  output [31:0] io_dout_bits,
  input         io_din_valid,
  input  [31:0] io_din_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] data; // @[util.scala 143:21]
  reg  valid; // @[util.scala 144:22]
  assign io_dout_valid = valid; // @[util.scala 151:17]
  assign io_dout_bits = data; // @[util.scala 152:16]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 143:21]
      data <= 32'h0; // @[util.scala 143:21]
    end else if (io_dout_ready) begin // @[util.scala 145:22]
      data <= io_din_bits; // @[util.scala 146:10]
    end
    if (reset) begin // @[util.scala 144:22]
      valid <= 1'h0; // @[util.scala 144:22]
    end else if (io_dout_ready) begin // @[util.scala 145:22]
      valid <= io_din_valid; // @[util.scala 147:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  valid = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pipeline_34(
  input        clock,
  input        reset,
  input        io_dout_ready,
  output       io_dout_valid,
  output [8:0] io_dout_bits,
  input        io_din_valid,
  input  [8:0] io_din_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] data; // @[util.scala 143:21]
  reg  valid; // @[util.scala 144:22]
  assign io_dout_valid = valid; // @[util.scala 151:17]
  assign io_dout_bits = data; // @[util.scala 152:16]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 143:21]
      data <= 9'h0; // @[util.scala 143:21]
    end else if (io_dout_ready) begin // @[util.scala 145:22]
      data <= io_din_bits; // @[util.scala 146:10]
    end
    if (reset) begin // @[util.scala 144:22]
      valid <= 1'h0; // @[util.scala 144:22]
    end else if (io_dout_ready) begin // @[util.scala 145:22]
      valid <= io_din_valid; // @[util.scala 147:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  valid = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h0; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_1(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h1; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_2(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h2; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_3(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h3; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_4(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h4; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_5(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h5; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_6(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h6; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_7(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h7; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_8(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h8; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_9(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'h9; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_10(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'ha; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_11(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'hb; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_12(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'hc; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_13(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'hd; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_14(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'he; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module Scatter_15(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata,
  output         io_end
);
  wire [16:0] bitmap__addra; // @[BFS.scala 705:22]
  wire  bitmap__clka; // @[BFS.scala 705:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 705:22]
  wire  bitmap__ena; // @[BFS.scala 705:22]
  wire  bitmap__wea; // @[BFS.scala 705:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 705:22]
  wire  bitmap__clkb; // @[BFS.scala 705:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 705:22]
  wire  bitmap__enb; // @[BFS.scala 705:22]
  wire  arbi_clock; // @[BFS.scala 706:20]
  wire  arbi_reset; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 706:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 706:20]
  wire [511:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 706:20]
  wire [15:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 706:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 706:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 706:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 739:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 739:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 739:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 739:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 740:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 740:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 740:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 740:31]
  wire  bitmap_wait_clock; // @[BFS.scala 749:27]
  wire  bitmap_wait_reset; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 749:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 749:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 749:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 754:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 754:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 759:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 759:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 759:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 764:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 764:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 764:41]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[3:0] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[35:32] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[67:64] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[99:96] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[131:128] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[163:160] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[195:192] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[227:224] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[259:256] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[291:288] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[323:320] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[355:352] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[387:384] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[419:416] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[451:448] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[BFS.scala 727:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[483:480] == 4'hf; // @[BFS.scala 709:39]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_5; // @[BFS.scala 728:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[BFS.scala 727:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 733:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8}; // @[BFS.scala 733:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 748:38]
  wire  _bitmap_write_addr_io_din_valid_T_1 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff; // @[BFS.scala 719:40]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[6:4]}; // @[BFS.scala 721:69 BFS.scala 721:69]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = bitmap_wait_io_dout_bits[30:4] > 27'he7fff ? 4'h8 :
    _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 719:8]
  wire [26:0] _bitmap_doutb_T_5 = bitmap_wait_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE = {{3'd0}, bitmap_wait_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 713:8]
  wire [26:0] _bitmap_doutb_T_12 = bitmap_write_addr_io_dout_bits[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{3'd0}, bitmap_write_addr_io_dout_bits[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_doutb_T_14 = bitmap_write_addr_io_dout_bits[30:4] > 27'he7fff ? _bitmap_doutb_T_12 :
    _bitmap_doutb_WIRE_1; // @[BFS.scala 713:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 771:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 770:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 756:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 756:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 762:61]
  wire [23:0] _GEN_0 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 762:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_0 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 762:49]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = vertex_in_fifo_dout[30:4] - 27'he7fff; // @[BFS.scala 714:38]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{3'd0}, vertex_in_fifo_dout[30:7]}; // @[BFS.scala 715:50 BFS.scala 715:50]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = vertex_in_fifo_dout[30:4] > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 713:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 766:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 112:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 705:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 706:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 739:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 740:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 749:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 754:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 759:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 764:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 737:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 790:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 793:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 112:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 788:19]
  assign bitmap__clka = clock; // @[BFS.scala 786:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 787:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 784:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 785:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 779:19]
  assign bitmap__clkb = clock; // @[BFS.scala 780:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 778:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 735:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 734:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 733:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 777:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 775:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 776:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 781:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 741:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 742:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 783:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 782:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 789:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 743:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 744:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 752:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 750:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 751:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 758:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 755:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 757:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 763:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 760:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 762:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 768:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 765:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 767:41]
endmodule
module axis_arbitrator_17(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [127:0] io_xbar_in_bits_tdata,
  input  [3:0]   io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] data; // @[BFS.scala 237:21]
  reg [3:0] keep; // @[BFS.scala 238:21]
  wire  _T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 240:25]
  wire  _select_T_1 = |keep[0]; // @[BFS.scala 246:125]
  wire  _select_T_4 = |keep[1]; // @[BFS.scala 246:125]
  wire  _select_T_7 = |keep[2]; // @[BFS.scala 246:125]
  wire  _select_T_10 = |keep[3]; // @[BFS.scala 246:125]
  wire [6:0] _select_T_12 = _select_T_10 ? 7'h8 : 7'h0; // @[Mux.scala 98:16]
  wire [6:0] _select_T_13 = _select_T_7 ? 7'h4 : _select_T_12; // @[Mux.scala 98:16]
  wire [6:0] _select_T_14 = _select_T_4 ? 7'h2 : _select_T_13; // @[Mux.scala 98:16]
  wire [6:0] select = _select_T_1 ? 7'h1 : _select_T_14; // @[Mux.scala 98:16]
  wire [31:0] _io_ddr_out_bits_tdata_T_8 = select[0] ? data[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_9 = select[1] ? data[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_10 = select[2] ? data[95:64] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_11 = select[3] ? data[127:96] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_12 = _io_ddr_out_bits_tdata_T_8 | _io_ddr_out_bits_tdata_T_9; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_13 = _io_ddr_out_bits_tdata_T_12 | _io_ddr_out_bits_tdata_T_10; // @[Mux.scala 27:72]
  wire  next_keep_0 = select[0] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_1 = select[1] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_2 = select[2] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire  next_keep_3 = select[3] ? 1'h0 : 1'h1; // @[BFS.scala 257:28]
  wire [3:0] _keep_T = {next_keep_3,next_keep_2,next_keep_1,next_keep_0}; // @[BFS.scala 262:36]
  wire [3:0] _keep_T_1 = keep & _keep_T; // @[BFS.scala 262:18]
  assign io_xbar_in_ready = ~(|keep); // @[BFS.scala 243:23]
  assign io_ddr_out_valid = |select; // @[BFS.scala 247:33]
  assign io_ddr_out_bits_tdata = _io_ddr_out_bits_tdata_T_13 | _io_ddr_out_bits_tdata_T_11; // @[Mux.scala 27:72]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 237:21]
      data <= 128'h0; // @[BFS.scala 237:21]
    end else if (io_xbar_in_valid & io_xbar_in_ready) begin // @[BFS.scala 240:45]
      data <= io_xbar_in_bits_tdata; // @[BFS.scala 241:10]
    end
    if (reset) begin // @[BFS.scala 238:21]
      keep <= 4'h0; // @[BFS.scala 238:21]
    end else if (_T) begin // @[BFS.scala 259:45]
      keep <= io_xbar_in_bits_tkeep; // @[BFS.scala 260:10]
    end else if (io_ddr_out_valid & io_ddr_out_ready) begin // @[BFS.scala 261:52]
      keep <= _keep_T_1; // @[BFS.scala 262:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  data = _RAND_0[127:0];
  _RAND_1 = {1{`RANDOM}};
  keep = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Gather(
  input          clock,
  input          reset,
  output         io_ddr_in_ready,
  input          io_ddr_in_valid,
  input  [511:0] io_ddr_in_bits_tdata,
  input  [15:0]  io_ddr_in_bits_tkeep,
  input          io_gather_out_0_ready,
  output         io_gather_out_0_valid,
  output [31:0]  io_gather_out_0_bits_tdata,
  input          io_gather_out_1_ready,
  output         io_gather_out_1_valid,
  output [31:0]  io_gather_out_1_bits_tdata,
  input          io_gather_out_2_ready,
  output         io_gather_out_2_valid,
  output [31:0]  io_gather_out_2_bits_tdata,
  input          io_gather_out_3_ready,
  output         io_gather_out_3_valid,
  output [31:0]  io_gather_out_3_bits_tdata,
  input          io_gather_out_4_ready,
  output         io_gather_out_4_valid,
  output [31:0]  io_gather_out_4_bits_tdata
);
  wire  broadcaster_aclk; // @[BFS.scala 274:27]
  wire  broadcaster_aresetn; // @[BFS.scala 274:27]
  wire [511:0] broadcaster_s_axis_tdata; // @[BFS.scala 274:27]
  wire [63:0] broadcaster_s_axis_tkeep; // @[BFS.scala 274:27]
  wire  broadcaster_s_axis_tlast; // @[BFS.scala 274:27]
  wire  broadcaster_s_axis_tvalid; // @[BFS.scala 274:27]
  wire  broadcaster_s_axis_tready; // @[BFS.scala 274:27]
  wire  broadcaster_s_axis_tid; // @[BFS.scala 274:27]
  wire [2559:0] broadcaster_m_axis_tdata; // @[BFS.scala 274:27]
  wire [319:0] broadcaster_m_axis_tkeep; // @[BFS.scala 274:27]
  wire [4:0] broadcaster_m_axis_tlast; // @[BFS.scala 274:27]
  wire [4:0] broadcaster_m_axis_tvalid; // @[BFS.scala 274:27]
  wire [4:0] broadcaster_m_axis_tready; // @[BFS.scala 274:27]
  wire [4:0] broadcaster_m_axis_tid; // @[BFS.scala 274:27]
  wire  v2Apply_fifo_s_axis_aclk; // @[BFS.scala 281:28]
  wire  v2Apply_fifo_s_axis_aresetn; // @[BFS.scala 281:28]
  wire [511:0] v2Apply_fifo_s_axis_tdata; // @[BFS.scala 281:28]
  wire [63:0] v2Apply_fifo_s_axis_tkeep; // @[BFS.scala 281:28]
  wire  v2Apply_fifo_s_axis_tlast; // @[BFS.scala 281:28]
  wire  v2Apply_fifo_s_axis_tvalid; // @[BFS.scala 281:28]
  wire  v2Apply_fifo_s_axis_tready; // @[BFS.scala 281:28]
  wire  v2Apply_fifo_s_axis_tid; // @[BFS.scala 281:28]
  wire [511:0] v2Apply_fifo_m_axis_tdata; // @[BFS.scala 281:28]
  wire [63:0] v2Apply_fifo_m_axis_tkeep; // @[BFS.scala 281:28]
  wire  v2Apply_fifo_m_axis_tlast; // @[BFS.scala 281:28]
  wire  v2Apply_fifo_m_axis_tvalid; // @[BFS.scala 281:28]
  wire  v2Apply_fifo_m_axis_tready; // @[BFS.scala 281:28]
  wire  v2Apply_fifo_m_axis_tid; // @[BFS.scala 281:28]
  wire  v2Broadcast_fifo_0_s_axis_aclk; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_0_s_axis_aresetn; // @[BFS.scala 290:16]
  wire [127:0] v2Broadcast_fifo_0_s_axis_tdata; // @[BFS.scala 290:16]
  wire [15:0] v2Broadcast_fifo_0_s_axis_tkeep; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_0_s_axis_tlast; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_0_s_axis_tvalid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_0_s_axis_tready; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_0_s_axis_tid; // @[BFS.scala 290:16]
  wire [127:0] v2Broadcast_fifo_0_m_axis_tdata; // @[BFS.scala 290:16]
  wire [15:0] v2Broadcast_fifo_0_m_axis_tkeep; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_0_m_axis_tlast; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_0_m_axis_tvalid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_0_m_axis_tready; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_0_m_axis_tid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_s_axis_aclk; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_s_axis_aresetn; // @[BFS.scala 290:16]
  wire [127:0] v2Broadcast_fifo_1_s_axis_tdata; // @[BFS.scala 290:16]
  wire [15:0] v2Broadcast_fifo_1_s_axis_tkeep; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_s_axis_tlast; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_s_axis_tvalid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_s_axis_tready; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_s_axis_tid; // @[BFS.scala 290:16]
  wire [127:0] v2Broadcast_fifo_1_m_axis_tdata; // @[BFS.scala 290:16]
  wire [15:0] v2Broadcast_fifo_1_m_axis_tkeep; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_m_axis_tlast; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_m_axis_tvalid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_m_axis_tready; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_1_m_axis_tid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_s_axis_aclk; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_s_axis_aresetn; // @[BFS.scala 290:16]
  wire [127:0] v2Broadcast_fifo_2_s_axis_tdata; // @[BFS.scala 290:16]
  wire [15:0] v2Broadcast_fifo_2_s_axis_tkeep; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_s_axis_tlast; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_s_axis_tvalid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_s_axis_tready; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_s_axis_tid; // @[BFS.scala 290:16]
  wire [127:0] v2Broadcast_fifo_2_m_axis_tdata; // @[BFS.scala 290:16]
  wire [15:0] v2Broadcast_fifo_2_m_axis_tkeep; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_m_axis_tlast; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_m_axis_tvalid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_m_axis_tready; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_2_m_axis_tid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_s_axis_aclk; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_s_axis_aresetn; // @[BFS.scala 290:16]
  wire [127:0] v2Broadcast_fifo_3_s_axis_tdata; // @[BFS.scala 290:16]
  wire [15:0] v2Broadcast_fifo_3_s_axis_tkeep; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_s_axis_tlast; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_s_axis_tvalid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_s_axis_tready; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_s_axis_tid; // @[BFS.scala 290:16]
  wire [127:0] v2Broadcast_fifo_3_m_axis_tdata; // @[BFS.scala 290:16]
  wire [15:0] v2Broadcast_fifo_3_m_axis_tkeep; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_m_axis_tlast; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_m_axis_tvalid; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_m_axis_tready; // @[BFS.scala 290:16]
  wire  v2Broadcast_fifo_3_m_axis_tid; // @[BFS.scala 290:16]
  wire  v2Apply_selecter_clock; // @[BFS.scala 319:32]
  wire  v2Apply_selecter_reset; // @[BFS.scala 319:32]
  wire  v2Apply_selecter_io_xbar_in_ready; // @[BFS.scala 319:32]
  wire  v2Apply_selecter_io_xbar_in_valid; // @[BFS.scala 319:32]
  wire [511:0] v2Apply_selecter_io_xbar_in_bits_tdata; // @[BFS.scala 319:32]
  wire [15:0] v2Apply_selecter_io_xbar_in_bits_tkeep; // @[BFS.scala 319:32]
  wire  v2Apply_selecter_io_ddr_out_ready; // @[BFS.scala 319:32]
  wire  v2Apply_selecter_io_ddr_out_valid; // @[BFS.scala 319:32]
  wire [31:0] v2Apply_selecter_io_ddr_out_bits_tdata; // @[BFS.scala 319:32]
  wire  v2Broadcast_selecter_0_clock; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_0_reset; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_ready; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_valid; // @[BFS.scala 326:16]
  wire [127:0] v2Broadcast_selecter_0_io_xbar_in_bits_tdata; // @[BFS.scala 326:16]
  wire [3:0] v2Broadcast_selecter_0_io_xbar_in_bits_tkeep; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_0_io_ddr_out_ready; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_0_io_ddr_out_valid; // @[BFS.scala 326:16]
  wire [31:0] v2Broadcast_selecter_0_io_ddr_out_bits_tdata; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_1_clock; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_1_reset; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_ready; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_valid; // @[BFS.scala 326:16]
  wire [127:0] v2Broadcast_selecter_1_io_xbar_in_bits_tdata; // @[BFS.scala 326:16]
  wire [3:0] v2Broadcast_selecter_1_io_xbar_in_bits_tkeep; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_1_io_ddr_out_ready; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_1_io_ddr_out_valid; // @[BFS.scala 326:16]
  wire [31:0] v2Broadcast_selecter_1_io_ddr_out_bits_tdata; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_2_clock; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_2_reset; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_ready; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_valid; // @[BFS.scala 326:16]
  wire [127:0] v2Broadcast_selecter_2_io_xbar_in_bits_tdata; // @[BFS.scala 326:16]
  wire [3:0] v2Broadcast_selecter_2_io_xbar_in_bits_tkeep; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_2_io_ddr_out_ready; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_2_io_ddr_out_valid; // @[BFS.scala 326:16]
  wire [31:0] v2Broadcast_selecter_2_io_ddr_out_bits_tdata; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_3_clock; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_3_reset; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_ready; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_valid; // @[BFS.scala 326:16]
  wire [127:0] v2Broadcast_selecter_3_io_xbar_in_bits_tdata; // @[BFS.scala 326:16]
  wire [3:0] v2Broadcast_selecter_3_io_xbar_in_bits_tkeep; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_3_io_ddr_out_ready; // @[BFS.scala 326:16]
  wire  v2Broadcast_selecter_3_io_ddr_out_valid; // @[BFS.scala 326:16]
  wire [31:0] v2Broadcast_selecter_3_io_ddr_out_bits_tdata; // @[BFS.scala 326:16]
  wire [63:0] v2Broadcast_fifo_0_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[159:128],broadcaster_m_axis_tdata[31:0]}
    ; // @[BFS.scala 299:16]
  wire [63:0] v2Broadcast_fifo_0_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[415:384],broadcaster_m_axis_tdata[287:
    256]}; // @[BFS.scala 299:16]
  wire  _v2Broadcast_fifo_0_io_s_axis_tvalid_T_29 = broadcaster_m_axis_tkeep[0] | broadcaster_m_axis_tkeep[4] |
    broadcaster_m_axis_tkeep[8] | broadcaster_m_axis_tkeep[12]; // @[BFS.scala 309:17]
  wire [3:0] _v2Broadcast_fifo_0_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[12],broadcaster_m_axis_tkeep[8],
    broadcaster_m_axis_tkeep[4],broadcaster_m_axis_tkeep[0]}; // @[BFS.scala 312:16]
  wire [63:0] v2Broadcast_fifo_1_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[703:672],broadcaster_m_axis_tdata[575:
    544]}; // @[BFS.scala 299:16]
  wire [63:0] v2Broadcast_fifo_1_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[959:928],broadcaster_m_axis_tdata[831:
    800]}; // @[BFS.scala 299:16]
  wire  _v2Broadcast_fifo_1_io_s_axis_tvalid_T_30 = broadcaster_m_axis_tkeep[1] | broadcaster_m_axis_tkeep[5] |
    broadcaster_m_axis_tkeep[9] | broadcaster_m_axis_tkeep[13]; // @[BFS.scala 309:17]
  wire [3:0] _v2Broadcast_fifo_1_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[13],broadcaster_m_axis_tkeep[9],
    broadcaster_m_axis_tkeep[5],broadcaster_m_axis_tkeep[1]}; // @[BFS.scala 312:16]
  wire [63:0] v2Broadcast_fifo_2_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[1247:1216],broadcaster_m_axis_tdata[1119
    :1088]}; // @[BFS.scala 299:16]
  wire [63:0] v2Broadcast_fifo_2_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[1503:1472],broadcaster_m_axis_tdata[1375
    :1344]}; // @[BFS.scala 299:16]
  wire  _v2Broadcast_fifo_2_io_s_axis_tvalid_T_31 = broadcaster_m_axis_tkeep[2] | broadcaster_m_axis_tkeep[6] |
    broadcaster_m_axis_tkeep[10] | broadcaster_m_axis_tkeep[14]; // @[BFS.scala 309:17]
  wire [3:0] _v2Broadcast_fifo_2_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[14],broadcaster_m_axis_tkeep[10],
    broadcaster_m_axis_tkeep[6],broadcaster_m_axis_tkeep[2]}; // @[BFS.scala 312:16]
  wire [63:0] v2Broadcast_fifo_3_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[1791:1760],broadcaster_m_axis_tdata[1663
    :1632]}; // @[BFS.scala 299:16]
  wire [63:0] v2Broadcast_fifo_3_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[2047:2016],broadcaster_m_axis_tdata[1919
    :1888]}; // @[BFS.scala 299:16]
  wire  _v2Broadcast_fifo_3_io_s_axis_tvalid_T_32 = broadcaster_m_axis_tkeep[3] | broadcaster_m_axis_tkeep[7] |
    broadcaster_m_axis_tkeep[11] | broadcaster_m_axis_tkeep[15]; // @[BFS.scala 309:17]
  wire [3:0] _v2Broadcast_fifo_3_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[15],broadcaster_m_axis_tkeep[11],
    broadcaster_m_axis_tkeep[7],broadcaster_m_axis_tkeep[3]}; // @[BFS.scala 312:16]
  wire  _broadcaster_io_m_axis_tready_WIRE_1 = v2Broadcast_fifo_1_s_axis_tready; // @[BFS.scala 317:101 BFS.scala 317:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_0 = v2Broadcast_fifo_0_s_axis_tready; // @[BFS.scala 317:101 BFS.scala 317:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_3 = v2Broadcast_fifo_3_s_axis_tready; // @[BFS.scala 317:101 BFS.scala 317:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_2 = v2Broadcast_fifo_2_s_axis_tready; // @[BFS.scala 317:101 BFS.scala 317:101]
  wire [3:0] broadcaster_io_m_axis_tready_lo_1 = {_broadcaster_io_m_axis_tready_WIRE_3,
    _broadcaster_io_m_axis_tready_WIRE_2,_broadcaster_io_m_axis_tready_WIRE_1,_broadcaster_io_m_axis_tready_WIRE_0}; // @[BFS.scala 317:151]
  wire [63:0] _v2Apply_selecter_io_xbar_in_bits_tkeep_T = v2Apply_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 113:21]
  wire [15:0] _v2Broadcast_selecter_0_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_0_m_axis_tkeep; // @[nf_arm_doce_top.scala 113:21]
  wire [15:0] _v2Broadcast_selecter_1_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_1_m_axis_tkeep; // @[nf_arm_doce_top.scala 113:21]
  wire [15:0] _v2Broadcast_selecter_2_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_2_m_axis_tkeep; // @[nf_arm_doce_top.scala 113:21]
  wire [15:0] _v2Broadcast_selecter_3_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_3_m_axis_tkeep; // @[nf_arm_doce_top.scala 113:21]
  gather_broadcaster broadcaster ( // @[BFS.scala 274:27]
    .aclk(broadcaster_aclk),
    .aresetn(broadcaster_aresetn),
    .s_axis_tdata(broadcaster_s_axis_tdata),
    .s_axis_tkeep(broadcaster_s_axis_tkeep),
    .s_axis_tlast(broadcaster_s_axis_tlast),
    .s_axis_tvalid(broadcaster_s_axis_tvalid),
    .s_axis_tready(broadcaster_s_axis_tready),
    .s_axis_tid(broadcaster_s_axis_tid),
    .m_axis_tdata(broadcaster_m_axis_tdata),
    .m_axis_tkeep(broadcaster_m_axis_tkeep),
    .m_axis_tlast(broadcaster_m_axis_tlast),
    .m_axis_tvalid(broadcaster_m_axis_tvalid),
    .m_axis_tready(broadcaster_m_axis_tready),
    .m_axis_tid(broadcaster_m_axis_tid)
  );
  v2A_fifo v2Apply_fifo ( // @[BFS.scala 281:28]
    .s_axis_aclk(v2Apply_fifo_s_axis_aclk),
    .s_axis_aresetn(v2Apply_fifo_s_axis_aresetn),
    .s_axis_tdata(v2Apply_fifo_s_axis_tdata),
    .s_axis_tkeep(v2Apply_fifo_s_axis_tkeep),
    .s_axis_tlast(v2Apply_fifo_s_axis_tlast),
    .s_axis_tvalid(v2Apply_fifo_s_axis_tvalid),
    .s_axis_tready(v2Apply_fifo_s_axis_tready),
    .s_axis_tid(v2Apply_fifo_s_axis_tid),
    .m_axis_tdata(v2Apply_fifo_m_axis_tdata),
    .m_axis_tkeep(v2Apply_fifo_m_axis_tkeep),
    .m_axis_tlast(v2Apply_fifo_m_axis_tlast),
    .m_axis_tvalid(v2Apply_fifo_m_axis_tvalid),
    .m_axis_tready(v2Apply_fifo_m_axis_tready),
    .m_axis_tid(v2Apply_fifo_m_axis_tid)
  );
  v2B_fifo v2Broadcast_fifo_0 ( // @[BFS.scala 290:16]
    .s_axis_aclk(v2Broadcast_fifo_0_s_axis_aclk),
    .s_axis_aresetn(v2Broadcast_fifo_0_s_axis_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_0_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_0_s_axis_tkeep),
    .s_axis_tlast(v2Broadcast_fifo_0_s_axis_tlast),
    .s_axis_tvalid(v2Broadcast_fifo_0_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_0_s_axis_tready),
    .s_axis_tid(v2Broadcast_fifo_0_s_axis_tid),
    .m_axis_tdata(v2Broadcast_fifo_0_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_0_m_axis_tkeep),
    .m_axis_tlast(v2Broadcast_fifo_0_m_axis_tlast),
    .m_axis_tvalid(v2Broadcast_fifo_0_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_0_m_axis_tready),
    .m_axis_tid(v2Broadcast_fifo_0_m_axis_tid)
  );
  v2B_fifo v2Broadcast_fifo_1 ( // @[BFS.scala 290:16]
    .s_axis_aclk(v2Broadcast_fifo_1_s_axis_aclk),
    .s_axis_aresetn(v2Broadcast_fifo_1_s_axis_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_1_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_1_s_axis_tkeep),
    .s_axis_tlast(v2Broadcast_fifo_1_s_axis_tlast),
    .s_axis_tvalid(v2Broadcast_fifo_1_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_1_s_axis_tready),
    .s_axis_tid(v2Broadcast_fifo_1_s_axis_tid),
    .m_axis_tdata(v2Broadcast_fifo_1_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_1_m_axis_tkeep),
    .m_axis_tlast(v2Broadcast_fifo_1_m_axis_tlast),
    .m_axis_tvalid(v2Broadcast_fifo_1_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_1_m_axis_tready),
    .m_axis_tid(v2Broadcast_fifo_1_m_axis_tid)
  );
  v2B_fifo v2Broadcast_fifo_2 ( // @[BFS.scala 290:16]
    .s_axis_aclk(v2Broadcast_fifo_2_s_axis_aclk),
    .s_axis_aresetn(v2Broadcast_fifo_2_s_axis_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_2_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_2_s_axis_tkeep),
    .s_axis_tlast(v2Broadcast_fifo_2_s_axis_tlast),
    .s_axis_tvalid(v2Broadcast_fifo_2_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_2_s_axis_tready),
    .s_axis_tid(v2Broadcast_fifo_2_s_axis_tid),
    .m_axis_tdata(v2Broadcast_fifo_2_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_2_m_axis_tkeep),
    .m_axis_tlast(v2Broadcast_fifo_2_m_axis_tlast),
    .m_axis_tvalid(v2Broadcast_fifo_2_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_2_m_axis_tready),
    .m_axis_tid(v2Broadcast_fifo_2_m_axis_tid)
  );
  v2B_fifo v2Broadcast_fifo_3 ( // @[BFS.scala 290:16]
    .s_axis_aclk(v2Broadcast_fifo_3_s_axis_aclk),
    .s_axis_aresetn(v2Broadcast_fifo_3_s_axis_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_3_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_3_s_axis_tkeep),
    .s_axis_tlast(v2Broadcast_fifo_3_s_axis_tlast),
    .s_axis_tvalid(v2Broadcast_fifo_3_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_3_s_axis_tready),
    .s_axis_tid(v2Broadcast_fifo_3_s_axis_tid),
    .m_axis_tdata(v2Broadcast_fifo_3_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_3_m_axis_tkeep),
    .m_axis_tlast(v2Broadcast_fifo_3_m_axis_tlast),
    .m_axis_tvalid(v2Broadcast_fifo_3_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_3_m_axis_tready),
    .m_axis_tid(v2Broadcast_fifo_3_m_axis_tid)
  );
  axis_arbitrator v2Apply_selecter ( // @[BFS.scala 319:32]
    .clock(v2Apply_selecter_clock),
    .reset(v2Apply_selecter_reset),
    .io_xbar_in_ready(v2Apply_selecter_io_xbar_in_ready),
    .io_xbar_in_valid(v2Apply_selecter_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Apply_selecter_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Apply_selecter_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Apply_selecter_io_ddr_out_ready),
    .io_ddr_out_valid(v2Apply_selecter_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Apply_selecter_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_17 v2Broadcast_selecter_0 ( // @[BFS.scala 326:16]
    .clock(v2Broadcast_selecter_0_clock),
    .reset(v2Broadcast_selecter_0_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_0_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_0_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Broadcast_selecter_0_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_0_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_0_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_17 v2Broadcast_selecter_1 ( // @[BFS.scala 326:16]
    .clock(v2Broadcast_selecter_1_clock),
    .reset(v2Broadcast_selecter_1_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_1_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_1_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Broadcast_selecter_1_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_1_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_1_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_17 v2Broadcast_selecter_2 ( // @[BFS.scala 326:16]
    .clock(v2Broadcast_selecter_2_clock),
    .reset(v2Broadcast_selecter_2_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_2_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_2_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Broadcast_selecter_2_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_2_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_2_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_17 v2Broadcast_selecter_3 ( // @[BFS.scala 326:16]
    .clock(v2Broadcast_selecter_3_clock),
    .reset(v2Broadcast_selecter_3_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_3_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_3_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Broadcast_selecter_3_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_3_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_3_io_ddr_out_bits_tdata)
  );
  assign io_ddr_in_ready = broadcaster_s_axis_tready; // @[BFS.scala 277:19]
  assign io_gather_out_0_valid = v2Broadcast_selecter_0_io_ddr_out_valid; // @[BFS.scala 333:20]
  assign io_gather_out_0_bits_tdata = v2Broadcast_selecter_0_io_ddr_out_bits_tdata; // @[BFS.scala 333:20]
  assign io_gather_out_1_valid = v2Broadcast_selecter_1_io_ddr_out_valid; // @[BFS.scala 333:20]
  assign io_gather_out_1_bits_tdata = v2Broadcast_selecter_1_io_ddr_out_bits_tdata; // @[BFS.scala 333:20]
  assign io_gather_out_2_valid = v2Broadcast_selecter_2_io_ddr_out_valid; // @[BFS.scala 333:20]
  assign io_gather_out_2_bits_tdata = v2Broadcast_selecter_2_io_ddr_out_bits_tdata; // @[BFS.scala 333:20]
  assign io_gather_out_3_valid = v2Broadcast_selecter_3_io_ddr_out_valid; // @[BFS.scala 333:20]
  assign io_gather_out_3_bits_tdata = v2Broadcast_selecter_3_io_ddr_out_bits_tdata; // @[BFS.scala 333:20]
  assign io_gather_out_4_valid = v2Apply_selecter_io_ddr_out_valid; // @[BFS.scala 323:31]
  assign io_gather_out_4_bits_tdata = v2Apply_selecter_io_ddr_out_bits_tdata; // @[BFS.scala 323:31]
  assign broadcaster_aclk = clock; // @[BFS.scala 279:38]
  assign broadcaster_aresetn = ~reset; // @[BFS.scala 278:29]
  assign broadcaster_s_axis_tdata = io_ddr_in_bits_tdata; // @[nf_arm_doce_top.scala 105:11]
  assign broadcaster_s_axis_tkeep = {{48'd0}, io_ddr_in_bits_tkeep}; // @[nf_arm_doce_top.scala 107:11]
  assign broadcaster_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 106:11]
  assign broadcaster_s_axis_tvalid = io_ddr_in_valid; // @[BFS.scala 276:32]
  assign broadcaster_s_axis_tid = 1'h0;
  assign broadcaster_m_axis_tready = {v2Apply_fifo_s_axis_tready,broadcaster_io_m_axis_tready_lo_1}; // @[Cat.scala 30:58]
  assign v2Apply_fifo_s_axis_aclk = clock; // @[BFS.scala 282:46]
  assign v2Apply_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 283:37]
  assign v2Apply_fifo_s_axis_tdata = broadcaster_m_axis_tdata[2559:2048]; // @[BFS.scala 284:62]
  assign v2Apply_fifo_s_axis_tkeep = broadcaster_m_axis_tkeep[319:256]; // @[BFS.scala 286:62]
  assign v2Apply_fifo_s_axis_tlast = broadcaster_m_axis_tlast[4]; // @[BFS.scala 287:62]
  assign v2Apply_fifo_s_axis_tvalid = broadcaster_m_axis_tvalid[4]; // @[BFS.scala 285:64]
  assign v2Apply_fifo_s_axis_tid = 1'h0;
  assign v2Apply_fifo_m_axis_tready = v2Apply_selecter_io_xbar_in_ready; // @[BFS.scala 321:33]
  assign v2Broadcast_fifo_0_s_axis_aclk = clock; // @[BFS.scala 295:39]
  assign v2Broadcast_fifo_0_s_axis_aresetn = ~reset; // @[BFS.scala 294:30]
  assign v2Broadcast_fifo_0_s_axis_tdata = {v2Broadcast_fifo_0_io_s_axis_tdata_hi,v2Broadcast_fifo_0_io_s_axis_tdata_lo}
    ; // @[BFS.scala 299:16]
  assign v2Broadcast_fifo_0_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_0_io_s_axis_tkeep_T_9}; // @[BFS.scala 312:16]
  assign v2Broadcast_fifo_0_s_axis_tlast = broadcaster_m_axis_tlast[0]; // @[BFS.scala 313:55]
  assign v2Broadcast_fifo_0_s_axis_tvalid = broadcaster_m_axis_tvalid[0] & _v2Broadcast_fifo_0_io_s_axis_tvalid_T_29; // @[BFS.scala 300:61]
  assign v2Broadcast_fifo_0_s_axis_tid = 1'h0;
  assign v2Broadcast_fifo_0_m_axis_tready = v2Broadcast_selecter_0_io_xbar_in_ready; // @[BFS.scala 332:44]
  assign v2Broadcast_fifo_1_s_axis_aclk = clock; // @[BFS.scala 295:39]
  assign v2Broadcast_fifo_1_s_axis_aresetn = ~reset; // @[BFS.scala 294:30]
  assign v2Broadcast_fifo_1_s_axis_tdata = {v2Broadcast_fifo_1_io_s_axis_tdata_hi,v2Broadcast_fifo_1_io_s_axis_tdata_lo}
    ; // @[BFS.scala 299:16]
  assign v2Broadcast_fifo_1_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_1_io_s_axis_tkeep_T_9}; // @[BFS.scala 312:16]
  assign v2Broadcast_fifo_1_s_axis_tlast = broadcaster_m_axis_tlast[1]; // @[BFS.scala 313:55]
  assign v2Broadcast_fifo_1_s_axis_tvalid = broadcaster_m_axis_tvalid[1] & _v2Broadcast_fifo_1_io_s_axis_tvalid_T_30; // @[BFS.scala 300:61]
  assign v2Broadcast_fifo_1_s_axis_tid = 1'h0;
  assign v2Broadcast_fifo_1_m_axis_tready = v2Broadcast_selecter_1_io_xbar_in_ready; // @[BFS.scala 332:44]
  assign v2Broadcast_fifo_2_s_axis_aclk = clock; // @[BFS.scala 295:39]
  assign v2Broadcast_fifo_2_s_axis_aresetn = ~reset; // @[BFS.scala 294:30]
  assign v2Broadcast_fifo_2_s_axis_tdata = {v2Broadcast_fifo_2_io_s_axis_tdata_hi,v2Broadcast_fifo_2_io_s_axis_tdata_lo}
    ; // @[BFS.scala 299:16]
  assign v2Broadcast_fifo_2_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_2_io_s_axis_tkeep_T_9}; // @[BFS.scala 312:16]
  assign v2Broadcast_fifo_2_s_axis_tlast = broadcaster_m_axis_tlast[2]; // @[BFS.scala 313:55]
  assign v2Broadcast_fifo_2_s_axis_tvalid = broadcaster_m_axis_tvalid[2] & _v2Broadcast_fifo_2_io_s_axis_tvalid_T_31; // @[BFS.scala 300:61]
  assign v2Broadcast_fifo_2_s_axis_tid = 1'h0;
  assign v2Broadcast_fifo_2_m_axis_tready = v2Broadcast_selecter_2_io_xbar_in_ready; // @[BFS.scala 332:44]
  assign v2Broadcast_fifo_3_s_axis_aclk = clock; // @[BFS.scala 295:39]
  assign v2Broadcast_fifo_3_s_axis_aresetn = ~reset; // @[BFS.scala 294:30]
  assign v2Broadcast_fifo_3_s_axis_tdata = {v2Broadcast_fifo_3_io_s_axis_tdata_hi,v2Broadcast_fifo_3_io_s_axis_tdata_lo}
    ; // @[BFS.scala 299:16]
  assign v2Broadcast_fifo_3_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_3_io_s_axis_tkeep_T_9}; // @[BFS.scala 312:16]
  assign v2Broadcast_fifo_3_s_axis_tlast = broadcaster_m_axis_tlast[3]; // @[BFS.scala 313:55]
  assign v2Broadcast_fifo_3_s_axis_tvalid = broadcaster_m_axis_tvalid[3] & _v2Broadcast_fifo_3_io_s_axis_tvalid_T_32; // @[BFS.scala 300:61]
  assign v2Broadcast_fifo_3_s_axis_tid = 1'h0;
  assign v2Broadcast_fifo_3_m_axis_tready = v2Broadcast_selecter_3_io_xbar_in_ready; // @[BFS.scala 332:44]
  assign v2Apply_selecter_clock = clock;
  assign v2Apply_selecter_reset = reset;
  assign v2Apply_selecter_io_xbar_in_valid = v2Apply_fifo_m_axis_tvalid; // @[BFS.scala 320:37]
  assign v2Apply_selecter_io_xbar_in_bits_tdata = v2Apply_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 111:21]
  assign v2Apply_selecter_io_xbar_in_bits_tkeep = _v2Apply_selecter_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 113:13]
  assign v2Apply_selecter_io_ddr_out_ready = io_gather_out_4_ready; // @[BFS.scala 323:31]
  assign v2Broadcast_selecter_0_clock = clock;
  assign v2Broadcast_selecter_0_reset = reset;
  assign v2Broadcast_selecter_0_io_xbar_in_valid = v2Broadcast_fifo_0_m_axis_tvalid; // @[BFS.scala 330:26]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tdata = v2Broadcast_fifo_0_m_axis_tdata; // @[nf_arm_doce_top.scala 111:21]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_0_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 113:13]
  assign v2Broadcast_selecter_0_io_ddr_out_ready = io_gather_out_0_ready; // @[BFS.scala 333:20]
  assign v2Broadcast_selecter_1_clock = clock;
  assign v2Broadcast_selecter_1_reset = reset;
  assign v2Broadcast_selecter_1_io_xbar_in_valid = v2Broadcast_fifo_1_m_axis_tvalid; // @[BFS.scala 330:26]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tdata = v2Broadcast_fifo_1_m_axis_tdata; // @[nf_arm_doce_top.scala 111:21]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_1_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 113:13]
  assign v2Broadcast_selecter_1_io_ddr_out_ready = io_gather_out_1_ready; // @[BFS.scala 333:20]
  assign v2Broadcast_selecter_2_clock = clock;
  assign v2Broadcast_selecter_2_reset = reset;
  assign v2Broadcast_selecter_2_io_xbar_in_valid = v2Broadcast_fifo_2_m_axis_tvalid; // @[BFS.scala 330:26]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tdata = v2Broadcast_fifo_2_m_axis_tdata; // @[nf_arm_doce_top.scala 111:21]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_2_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 113:13]
  assign v2Broadcast_selecter_2_io_ddr_out_ready = io_gather_out_2_ready; // @[BFS.scala 333:20]
  assign v2Broadcast_selecter_3_clock = clock;
  assign v2Broadcast_selecter_3_reset = reset;
  assign v2Broadcast_selecter_3_io_xbar_in_valid = v2Broadcast_fifo_3_m_axis_tvalid; // @[BFS.scala 330:26]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tdata = v2Broadcast_fifo_3_m_axis_tdata; // @[nf_arm_doce_top.scala 111:21]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_3_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 113:13]
  assign v2Broadcast_selecter_3_io_ddr_out_ready = io_gather_out_3_ready; // @[BFS.scala 333:20]
endmodule
module URAM_cluster(
  input  [17:0] io_addra,
  input         io_clka,
  input  [47:0] io_dina,
  input         io_wea,
  input  [17:0] io_addrb,
  input         io_clkb,
  output [47:0] io_doutb
);
  wire [11:0] cluster_0_addra; // @[util.scala 28:45]
  wire  cluster_0_clka; // @[util.scala 28:45]
  wire [47:0] cluster_0_dina; // @[util.scala 28:45]
  wire [47:0] cluster_0_douta; // @[util.scala 28:45]
  wire  cluster_0_ena; // @[util.scala 28:45]
  wire  cluster_0_wea; // @[util.scala 28:45]
  wire [11:0] cluster_0_addrb; // @[util.scala 28:45]
  wire  cluster_0_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_0_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_0_doutb; // @[util.scala 28:45]
  wire  cluster_0_enb; // @[util.scala 28:45]
  wire  cluster_0_web; // @[util.scala 28:45]
  wire [11:0] cluster_1_addra; // @[util.scala 28:45]
  wire  cluster_1_clka; // @[util.scala 28:45]
  wire [47:0] cluster_1_dina; // @[util.scala 28:45]
  wire [47:0] cluster_1_douta; // @[util.scala 28:45]
  wire  cluster_1_ena; // @[util.scala 28:45]
  wire  cluster_1_wea; // @[util.scala 28:45]
  wire [11:0] cluster_1_addrb; // @[util.scala 28:45]
  wire  cluster_1_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_1_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_1_doutb; // @[util.scala 28:45]
  wire  cluster_1_enb; // @[util.scala 28:45]
  wire  cluster_1_web; // @[util.scala 28:45]
  wire [11:0] cluster_2_addra; // @[util.scala 28:45]
  wire  cluster_2_clka; // @[util.scala 28:45]
  wire [47:0] cluster_2_dina; // @[util.scala 28:45]
  wire [47:0] cluster_2_douta; // @[util.scala 28:45]
  wire  cluster_2_ena; // @[util.scala 28:45]
  wire  cluster_2_wea; // @[util.scala 28:45]
  wire [11:0] cluster_2_addrb; // @[util.scala 28:45]
  wire  cluster_2_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_2_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_2_doutb; // @[util.scala 28:45]
  wire  cluster_2_enb; // @[util.scala 28:45]
  wire  cluster_2_web; // @[util.scala 28:45]
  wire [11:0] cluster_3_addra; // @[util.scala 28:45]
  wire  cluster_3_clka; // @[util.scala 28:45]
  wire [47:0] cluster_3_dina; // @[util.scala 28:45]
  wire [47:0] cluster_3_douta; // @[util.scala 28:45]
  wire  cluster_3_ena; // @[util.scala 28:45]
  wire  cluster_3_wea; // @[util.scala 28:45]
  wire [11:0] cluster_3_addrb; // @[util.scala 28:45]
  wire  cluster_3_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_3_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_3_doutb; // @[util.scala 28:45]
  wire  cluster_3_enb; // @[util.scala 28:45]
  wire  cluster_3_web; // @[util.scala 28:45]
  wire [11:0] cluster_4_addra; // @[util.scala 28:45]
  wire  cluster_4_clka; // @[util.scala 28:45]
  wire [47:0] cluster_4_dina; // @[util.scala 28:45]
  wire [47:0] cluster_4_douta; // @[util.scala 28:45]
  wire  cluster_4_ena; // @[util.scala 28:45]
  wire  cluster_4_wea; // @[util.scala 28:45]
  wire [11:0] cluster_4_addrb; // @[util.scala 28:45]
  wire  cluster_4_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_4_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_4_doutb; // @[util.scala 28:45]
  wire  cluster_4_enb; // @[util.scala 28:45]
  wire  cluster_4_web; // @[util.scala 28:45]
  wire [11:0] cluster_5_addra; // @[util.scala 28:45]
  wire  cluster_5_clka; // @[util.scala 28:45]
  wire [47:0] cluster_5_dina; // @[util.scala 28:45]
  wire [47:0] cluster_5_douta; // @[util.scala 28:45]
  wire  cluster_5_ena; // @[util.scala 28:45]
  wire  cluster_5_wea; // @[util.scala 28:45]
  wire [11:0] cluster_5_addrb; // @[util.scala 28:45]
  wire  cluster_5_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_5_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_5_doutb; // @[util.scala 28:45]
  wire  cluster_5_enb; // @[util.scala 28:45]
  wire  cluster_5_web; // @[util.scala 28:45]
  wire [11:0] cluster_6_addra; // @[util.scala 28:45]
  wire  cluster_6_clka; // @[util.scala 28:45]
  wire [47:0] cluster_6_dina; // @[util.scala 28:45]
  wire [47:0] cluster_6_douta; // @[util.scala 28:45]
  wire  cluster_6_ena; // @[util.scala 28:45]
  wire  cluster_6_wea; // @[util.scala 28:45]
  wire [11:0] cluster_6_addrb; // @[util.scala 28:45]
  wire  cluster_6_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_6_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_6_doutb; // @[util.scala 28:45]
  wire  cluster_6_enb; // @[util.scala 28:45]
  wire  cluster_6_web; // @[util.scala 28:45]
  wire [11:0] cluster_7_addra; // @[util.scala 28:45]
  wire  cluster_7_clka; // @[util.scala 28:45]
  wire [47:0] cluster_7_dina; // @[util.scala 28:45]
  wire [47:0] cluster_7_douta; // @[util.scala 28:45]
  wire  cluster_7_ena; // @[util.scala 28:45]
  wire  cluster_7_wea; // @[util.scala 28:45]
  wire [11:0] cluster_7_addrb; // @[util.scala 28:45]
  wire  cluster_7_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_7_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_7_doutb; // @[util.scala 28:45]
  wire  cluster_7_enb; // @[util.scala 28:45]
  wire  cluster_7_web; // @[util.scala 28:45]
  wire [11:0] cluster_8_addra; // @[util.scala 28:45]
  wire  cluster_8_clka; // @[util.scala 28:45]
  wire [47:0] cluster_8_dina; // @[util.scala 28:45]
  wire [47:0] cluster_8_douta; // @[util.scala 28:45]
  wire  cluster_8_ena; // @[util.scala 28:45]
  wire  cluster_8_wea; // @[util.scala 28:45]
  wire [11:0] cluster_8_addrb; // @[util.scala 28:45]
  wire  cluster_8_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_8_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_8_doutb; // @[util.scala 28:45]
  wire  cluster_8_enb; // @[util.scala 28:45]
  wire  cluster_8_web; // @[util.scala 28:45]
  wire [11:0] cluster_9_addra; // @[util.scala 28:45]
  wire  cluster_9_clka; // @[util.scala 28:45]
  wire [47:0] cluster_9_dina; // @[util.scala 28:45]
  wire [47:0] cluster_9_douta; // @[util.scala 28:45]
  wire  cluster_9_ena; // @[util.scala 28:45]
  wire  cluster_9_wea; // @[util.scala 28:45]
  wire [11:0] cluster_9_addrb; // @[util.scala 28:45]
  wire  cluster_9_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_9_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_9_doutb; // @[util.scala 28:45]
  wire  cluster_9_enb; // @[util.scala 28:45]
  wire  cluster_9_web; // @[util.scala 28:45]
  wire [11:0] cluster_10_addra; // @[util.scala 28:45]
  wire  cluster_10_clka; // @[util.scala 28:45]
  wire [47:0] cluster_10_dina; // @[util.scala 28:45]
  wire [47:0] cluster_10_douta; // @[util.scala 28:45]
  wire  cluster_10_ena; // @[util.scala 28:45]
  wire  cluster_10_wea; // @[util.scala 28:45]
  wire [11:0] cluster_10_addrb; // @[util.scala 28:45]
  wire  cluster_10_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_10_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_10_doutb; // @[util.scala 28:45]
  wire  cluster_10_enb; // @[util.scala 28:45]
  wire  cluster_10_web; // @[util.scala 28:45]
  wire [11:0] cluster_11_addra; // @[util.scala 28:45]
  wire  cluster_11_clka; // @[util.scala 28:45]
  wire [47:0] cluster_11_dina; // @[util.scala 28:45]
  wire [47:0] cluster_11_douta; // @[util.scala 28:45]
  wire  cluster_11_ena; // @[util.scala 28:45]
  wire  cluster_11_wea; // @[util.scala 28:45]
  wire [11:0] cluster_11_addrb; // @[util.scala 28:45]
  wire  cluster_11_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_11_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_11_doutb; // @[util.scala 28:45]
  wire  cluster_11_enb; // @[util.scala 28:45]
  wire  cluster_11_web; // @[util.scala 28:45]
  wire [11:0] cluster_12_addra; // @[util.scala 28:45]
  wire  cluster_12_clka; // @[util.scala 28:45]
  wire [47:0] cluster_12_dina; // @[util.scala 28:45]
  wire [47:0] cluster_12_douta; // @[util.scala 28:45]
  wire  cluster_12_ena; // @[util.scala 28:45]
  wire  cluster_12_wea; // @[util.scala 28:45]
  wire [11:0] cluster_12_addrb; // @[util.scala 28:45]
  wire  cluster_12_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_12_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_12_doutb; // @[util.scala 28:45]
  wire  cluster_12_enb; // @[util.scala 28:45]
  wire  cluster_12_web; // @[util.scala 28:45]
  wire [11:0] cluster_13_addra; // @[util.scala 28:45]
  wire  cluster_13_clka; // @[util.scala 28:45]
  wire [47:0] cluster_13_dina; // @[util.scala 28:45]
  wire [47:0] cluster_13_douta; // @[util.scala 28:45]
  wire  cluster_13_ena; // @[util.scala 28:45]
  wire  cluster_13_wea; // @[util.scala 28:45]
  wire [11:0] cluster_13_addrb; // @[util.scala 28:45]
  wire  cluster_13_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_13_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_13_doutb; // @[util.scala 28:45]
  wire  cluster_13_enb; // @[util.scala 28:45]
  wire  cluster_13_web; // @[util.scala 28:45]
  wire [11:0] cluster_14_addra; // @[util.scala 28:45]
  wire  cluster_14_clka; // @[util.scala 28:45]
  wire [47:0] cluster_14_dina; // @[util.scala 28:45]
  wire [47:0] cluster_14_douta; // @[util.scala 28:45]
  wire  cluster_14_ena; // @[util.scala 28:45]
  wire  cluster_14_wea; // @[util.scala 28:45]
  wire [11:0] cluster_14_addrb; // @[util.scala 28:45]
  wire  cluster_14_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_14_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_14_doutb; // @[util.scala 28:45]
  wire  cluster_14_enb; // @[util.scala 28:45]
  wire  cluster_14_web; // @[util.scala 28:45]
  wire [11:0] cluster_15_addra; // @[util.scala 28:45]
  wire  cluster_15_clka; // @[util.scala 28:45]
  wire [47:0] cluster_15_dina; // @[util.scala 28:45]
  wire [47:0] cluster_15_douta; // @[util.scala 28:45]
  wire  cluster_15_ena; // @[util.scala 28:45]
  wire  cluster_15_wea; // @[util.scala 28:45]
  wire [11:0] cluster_15_addrb; // @[util.scala 28:45]
  wire  cluster_15_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_15_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_15_doutb; // @[util.scala 28:45]
  wire  cluster_15_enb; // @[util.scala 28:45]
  wire  cluster_15_web; // @[util.scala 28:45]
  wire [11:0] cluster_16_addra; // @[util.scala 28:45]
  wire  cluster_16_clka; // @[util.scala 28:45]
  wire [47:0] cluster_16_dina; // @[util.scala 28:45]
  wire [47:0] cluster_16_douta; // @[util.scala 28:45]
  wire  cluster_16_ena; // @[util.scala 28:45]
  wire  cluster_16_wea; // @[util.scala 28:45]
  wire [11:0] cluster_16_addrb; // @[util.scala 28:45]
  wire  cluster_16_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_16_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_16_doutb; // @[util.scala 28:45]
  wire  cluster_16_enb; // @[util.scala 28:45]
  wire  cluster_16_web; // @[util.scala 28:45]
  wire [11:0] cluster_17_addra; // @[util.scala 28:45]
  wire  cluster_17_clka; // @[util.scala 28:45]
  wire [47:0] cluster_17_dina; // @[util.scala 28:45]
  wire [47:0] cluster_17_douta; // @[util.scala 28:45]
  wire  cluster_17_ena; // @[util.scala 28:45]
  wire  cluster_17_wea; // @[util.scala 28:45]
  wire [11:0] cluster_17_addrb; // @[util.scala 28:45]
  wire  cluster_17_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_17_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_17_doutb; // @[util.scala 28:45]
  wire  cluster_17_enb; // @[util.scala 28:45]
  wire  cluster_17_web; // @[util.scala 28:45]
  wire [11:0] cluster_18_addra; // @[util.scala 28:45]
  wire  cluster_18_clka; // @[util.scala 28:45]
  wire [47:0] cluster_18_dina; // @[util.scala 28:45]
  wire [47:0] cluster_18_douta; // @[util.scala 28:45]
  wire  cluster_18_ena; // @[util.scala 28:45]
  wire  cluster_18_wea; // @[util.scala 28:45]
  wire [11:0] cluster_18_addrb; // @[util.scala 28:45]
  wire  cluster_18_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_18_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_18_doutb; // @[util.scala 28:45]
  wire  cluster_18_enb; // @[util.scala 28:45]
  wire  cluster_18_web; // @[util.scala 28:45]
  wire [11:0] cluster_19_addra; // @[util.scala 28:45]
  wire  cluster_19_clka; // @[util.scala 28:45]
  wire [47:0] cluster_19_dina; // @[util.scala 28:45]
  wire [47:0] cluster_19_douta; // @[util.scala 28:45]
  wire  cluster_19_ena; // @[util.scala 28:45]
  wire  cluster_19_wea; // @[util.scala 28:45]
  wire [11:0] cluster_19_addrb; // @[util.scala 28:45]
  wire  cluster_19_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_19_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_19_doutb; // @[util.scala 28:45]
  wire  cluster_19_enb; // @[util.scala 28:45]
  wire  cluster_19_web; // @[util.scala 28:45]
  wire [11:0] cluster_20_addra; // @[util.scala 28:45]
  wire  cluster_20_clka; // @[util.scala 28:45]
  wire [47:0] cluster_20_dina; // @[util.scala 28:45]
  wire [47:0] cluster_20_douta; // @[util.scala 28:45]
  wire  cluster_20_ena; // @[util.scala 28:45]
  wire  cluster_20_wea; // @[util.scala 28:45]
  wire [11:0] cluster_20_addrb; // @[util.scala 28:45]
  wire  cluster_20_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_20_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_20_doutb; // @[util.scala 28:45]
  wire  cluster_20_enb; // @[util.scala 28:45]
  wire  cluster_20_web; // @[util.scala 28:45]
  wire [11:0] cluster_21_addra; // @[util.scala 28:45]
  wire  cluster_21_clka; // @[util.scala 28:45]
  wire [47:0] cluster_21_dina; // @[util.scala 28:45]
  wire [47:0] cluster_21_douta; // @[util.scala 28:45]
  wire  cluster_21_ena; // @[util.scala 28:45]
  wire  cluster_21_wea; // @[util.scala 28:45]
  wire [11:0] cluster_21_addrb; // @[util.scala 28:45]
  wire  cluster_21_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_21_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_21_doutb; // @[util.scala 28:45]
  wire  cluster_21_enb; // @[util.scala 28:45]
  wire  cluster_21_web; // @[util.scala 28:45]
  wire [11:0] cluster_22_addra; // @[util.scala 28:45]
  wire  cluster_22_clka; // @[util.scala 28:45]
  wire [47:0] cluster_22_dina; // @[util.scala 28:45]
  wire [47:0] cluster_22_douta; // @[util.scala 28:45]
  wire  cluster_22_ena; // @[util.scala 28:45]
  wire  cluster_22_wea; // @[util.scala 28:45]
  wire [11:0] cluster_22_addrb; // @[util.scala 28:45]
  wire  cluster_22_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_22_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_22_doutb; // @[util.scala 28:45]
  wire  cluster_22_enb; // @[util.scala 28:45]
  wire  cluster_22_web; // @[util.scala 28:45]
  wire [11:0] cluster_23_addra; // @[util.scala 28:45]
  wire  cluster_23_clka; // @[util.scala 28:45]
  wire [47:0] cluster_23_dina; // @[util.scala 28:45]
  wire [47:0] cluster_23_douta; // @[util.scala 28:45]
  wire  cluster_23_ena; // @[util.scala 28:45]
  wire  cluster_23_wea; // @[util.scala 28:45]
  wire [11:0] cluster_23_addrb; // @[util.scala 28:45]
  wire  cluster_23_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_23_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_23_doutb; // @[util.scala 28:45]
  wire  cluster_23_enb; // @[util.scala 28:45]
  wire  cluster_23_web; // @[util.scala 28:45]
  wire [11:0] cluster_24_addra; // @[util.scala 28:45]
  wire  cluster_24_clka; // @[util.scala 28:45]
  wire [47:0] cluster_24_dina; // @[util.scala 28:45]
  wire [47:0] cluster_24_douta; // @[util.scala 28:45]
  wire  cluster_24_ena; // @[util.scala 28:45]
  wire  cluster_24_wea; // @[util.scala 28:45]
  wire [11:0] cluster_24_addrb; // @[util.scala 28:45]
  wire  cluster_24_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_24_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_24_doutb; // @[util.scala 28:45]
  wire  cluster_24_enb; // @[util.scala 28:45]
  wire  cluster_24_web; // @[util.scala 28:45]
  wire [11:0] cluster_25_addra; // @[util.scala 28:45]
  wire  cluster_25_clka; // @[util.scala 28:45]
  wire [47:0] cluster_25_dina; // @[util.scala 28:45]
  wire [47:0] cluster_25_douta; // @[util.scala 28:45]
  wire  cluster_25_ena; // @[util.scala 28:45]
  wire  cluster_25_wea; // @[util.scala 28:45]
  wire [11:0] cluster_25_addrb; // @[util.scala 28:45]
  wire  cluster_25_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_25_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_25_doutb; // @[util.scala 28:45]
  wire  cluster_25_enb; // @[util.scala 28:45]
  wire  cluster_25_web; // @[util.scala 28:45]
  wire [11:0] cluster_26_addra; // @[util.scala 28:45]
  wire  cluster_26_clka; // @[util.scala 28:45]
  wire [47:0] cluster_26_dina; // @[util.scala 28:45]
  wire [47:0] cluster_26_douta; // @[util.scala 28:45]
  wire  cluster_26_ena; // @[util.scala 28:45]
  wire  cluster_26_wea; // @[util.scala 28:45]
  wire [11:0] cluster_26_addrb; // @[util.scala 28:45]
  wire  cluster_26_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_26_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_26_doutb; // @[util.scala 28:45]
  wire  cluster_26_enb; // @[util.scala 28:45]
  wire  cluster_26_web; // @[util.scala 28:45]
  wire [11:0] cluster_27_addra; // @[util.scala 28:45]
  wire  cluster_27_clka; // @[util.scala 28:45]
  wire [47:0] cluster_27_dina; // @[util.scala 28:45]
  wire [47:0] cluster_27_douta; // @[util.scala 28:45]
  wire  cluster_27_ena; // @[util.scala 28:45]
  wire  cluster_27_wea; // @[util.scala 28:45]
  wire [11:0] cluster_27_addrb; // @[util.scala 28:45]
  wire  cluster_27_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_27_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_27_doutb; // @[util.scala 28:45]
  wire  cluster_27_enb; // @[util.scala 28:45]
  wire  cluster_27_web; // @[util.scala 28:45]
  wire [11:0] cluster_28_addra; // @[util.scala 28:45]
  wire  cluster_28_clka; // @[util.scala 28:45]
  wire [47:0] cluster_28_dina; // @[util.scala 28:45]
  wire [47:0] cluster_28_douta; // @[util.scala 28:45]
  wire  cluster_28_ena; // @[util.scala 28:45]
  wire  cluster_28_wea; // @[util.scala 28:45]
  wire [11:0] cluster_28_addrb; // @[util.scala 28:45]
  wire  cluster_28_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_28_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_28_doutb; // @[util.scala 28:45]
  wire  cluster_28_enb; // @[util.scala 28:45]
  wire  cluster_28_web; // @[util.scala 28:45]
  wire [11:0] cluster_29_addra; // @[util.scala 28:45]
  wire  cluster_29_clka; // @[util.scala 28:45]
  wire [47:0] cluster_29_dina; // @[util.scala 28:45]
  wire [47:0] cluster_29_douta; // @[util.scala 28:45]
  wire  cluster_29_ena; // @[util.scala 28:45]
  wire  cluster_29_wea; // @[util.scala 28:45]
  wire [11:0] cluster_29_addrb; // @[util.scala 28:45]
  wire  cluster_29_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_29_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_29_doutb; // @[util.scala 28:45]
  wire  cluster_29_enb; // @[util.scala 28:45]
  wire  cluster_29_web; // @[util.scala 28:45]
  wire [11:0] cluster_30_addra; // @[util.scala 28:45]
  wire  cluster_30_clka; // @[util.scala 28:45]
  wire [47:0] cluster_30_dina; // @[util.scala 28:45]
  wire [47:0] cluster_30_douta; // @[util.scala 28:45]
  wire  cluster_30_ena; // @[util.scala 28:45]
  wire  cluster_30_wea; // @[util.scala 28:45]
  wire [11:0] cluster_30_addrb; // @[util.scala 28:45]
  wire  cluster_30_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_30_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_30_doutb; // @[util.scala 28:45]
  wire  cluster_30_enb; // @[util.scala 28:45]
  wire  cluster_30_web; // @[util.scala 28:45]
  wire [11:0] cluster_31_addra; // @[util.scala 28:45]
  wire  cluster_31_clka; // @[util.scala 28:45]
  wire [47:0] cluster_31_dina; // @[util.scala 28:45]
  wire [47:0] cluster_31_douta; // @[util.scala 28:45]
  wire  cluster_31_ena; // @[util.scala 28:45]
  wire  cluster_31_wea; // @[util.scala 28:45]
  wire [11:0] cluster_31_addrb; // @[util.scala 28:45]
  wire  cluster_31_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_31_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_31_doutb; // @[util.scala 28:45]
  wire  cluster_31_enb; // @[util.scala 28:45]
  wire  cluster_31_web; // @[util.scala 28:45]
  wire [11:0] cluster_32_addra; // @[util.scala 28:45]
  wire  cluster_32_clka; // @[util.scala 28:45]
  wire [47:0] cluster_32_dina; // @[util.scala 28:45]
  wire [47:0] cluster_32_douta; // @[util.scala 28:45]
  wire  cluster_32_ena; // @[util.scala 28:45]
  wire  cluster_32_wea; // @[util.scala 28:45]
  wire [11:0] cluster_32_addrb; // @[util.scala 28:45]
  wire  cluster_32_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_32_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_32_doutb; // @[util.scala 28:45]
  wire  cluster_32_enb; // @[util.scala 28:45]
  wire  cluster_32_web; // @[util.scala 28:45]
  wire [11:0] cluster_33_addra; // @[util.scala 28:45]
  wire  cluster_33_clka; // @[util.scala 28:45]
  wire [47:0] cluster_33_dina; // @[util.scala 28:45]
  wire [47:0] cluster_33_douta; // @[util.scala 28:45]
  wire  cluster_33_ena; // @[util.scala 28:45]
  wire  cluster_33_wea; // @[util.scala 28:45]
  wire [11:0] cluster_33_addrb; // @[util.scala 28:45]
  wire  cluster_33_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_33_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_33_doutb; // @[util.scala 28:45]
  wire  cluster_33_enb; // @[util.scala 28:45]
  wire  cluster_33_web; // @[util.scala 28:45]
  wire [11:0] cluster_34_addra; // @[util.scala 28:45]
  wire  cluster_34_clka; // @[util.scala 28:45]
  wire [47:0] cluster_34_dina; // @[util.scala 28:45]
  wire [47:0] cluster_34_douta; // @[util.scala 28:45]
  wire  cluster_34_ena; // @[util.scala 28:45]
  wire  cluster_34_wea; // @[util.scala 28:45]
  wire [11:0] cluster_34_addrb; // @[util.scala 28:45]
  wire  cluster_34_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_34_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_34_doutb; // @[util.scala 28:45]
  wire  cluster_34_enb; // @[util.scala 28:45]
  wire  cluster_34_web; // @[util.scala 28:45]
  wire [11:0] cluster_35_addra; // @[util.scala 28:45]
  wire  cluster_35_clka; // @[util.scala 28:45]
  wire [47:0] cluster_35_dina; // @[util.scala 28:45]
  wire [47:0] cluster_35_douta; // @[util.scala 28:45]
  wire  cluster_35_ena; // @[util.scala 28:45]
  wire  cluster_35_wea; // @[util.scala 28:45]
  wire [11:0] cluster_35_addrb; // @[util.scala 28:45]
  wire  cluster_35_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_35_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_35_doutb; // @[util.scala 28:45]
  wire  cluster_35_enb; // @[util.scala 28:45]
  wire  cluster_35_web; // @[util.scala 28:45]
  wire [11:0] cluster_36_addra; // @[util.scala 28:45]
  wire  cluster_36_clka; // @[util.scala 28:45]
  wire [47:0] cluster_36_dina; // @[util.scala 28:45]
  wire [47:0] cluster_36_douta; // @[util.scala 28:45]
  wire  cluster_36_ena; // @[util.scala 28:45]
  wire  cluster_36_wea; // @[util.scala 28:45]
  wire [11:0] cluster_36_addrb; // @[util.scala 28:45]
  wire  cluster_36_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_36_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_36_doutb; // @[util.scala 28:45]
  wire  cluster_36_enb; // @[util.scala 28:45]
  wire  cluster_36_web; // @[util.scala 28:45]
  wire [11:0] cluster_37_addra; // @[util.scala 28:45]
  wire  cluster_37_clka; // @[util.scala 28:45]
  wire [47:0] cluster_37_dina; // @[util.scala 28:45]
  wire [47:0] cluster_37_douta; // @[util.scala 28:45]
  wire  cluster_37_ena; // @[util.scala 28:45]
  wire  cluster_37_wea; // @[util.scala 28:45]
  wire [11:0] cluster_37_addrb; // @[util.scala 28:45]
  wire  cluster_37_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_37_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_37_doutb; // @[util.scala 28:45]
  wire  cluster_37_enb; // @[util.scala 28:45]
  wire  cluster_37_web; // @[util.scala 28:45]
  wire [11:0] cluster_38_addra; // @[util.scala 28:45]
  wire  cluster_38_clka; // @[util.scala 28:45]
  wire [47:0] cluster_38_dina; // @[util.scala 28:45]
  wire [47:0] cluster_38_douta; // @[util.scala 28:45]
  wire  cluster_38_ena; // @[util.scala 28:45]
  wire  cluster_38_wea; // @[util.scala 28:45]
  wire [11:0] cluster_38_addrb; // @[util.scala 28:45]
  wire  cluster_38_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_38_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_38_doutb; // @[util.scala 28:45]
  wire  cluster_38_enb; // @[util.scala 28:45]
  wire  cluster_38_web; // @[util.scala 28:45]
  wire [11:0] cluster_39_addra; // @[util.scala 28:45]
  wire  cluster_39_clka; // @[util.scala 28:45]
  wire [47:0] cluster_39_dina; // @[util.scala 28:45]
  wire [47:0] cluster_39_douta; // @[util.scala 28:45]
  wire  cluster_39_ena; // @[util.scala 28:45]
  wire  cluster_39_wea; // @[util.scala 28:45]
  wire [11:0] cluster_39_addrb; // @[util.scala 28:45]
  wire  cluster_39_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_39_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_39_doutb; // @[util.scala 28:45]
  wire  cluster_39_enb; // @[util.scala 28:45]
  wire  cluster_39_web; // @[util.scala 28:45]
  wire [11:0] cluster_40_addra; // @[util.scala 28:45]
  wire  cluster_40_clka; // @[util.scala 28:45]
  wire [47:0] cluster_40_dina; // @[util.scala 28:45]
  wire [47:0] cluster_40_douta; // @[util.scala 28:45]
  wire  cluster_40_ena; // @[util.scala 28:45]
  wire  cluster_40_wea; // @[util.scala 28:45]
  wire [11:0] cluster_40_addrb; // @[util.scala 28:45]
  wire  cluster_40_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_40_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_40_doutb; // @[util.scala 28:45]
  wire  cluster_40_enb; // @[util.scala 28:45]
  wire  cluster_40_web; // @[util.scala 28:45]
  wire [11:0] cluster_41_addra; // @[util.scala 28:45]
  wire  cluster_41_clka; // @[util.scala 28:45]
  wire [47:0] cluster_41_dina; // @[util.scala 28:45]
  wire [47:0] cluster_41_douta; // @[util.scala 28:45]
  wire  cluster_41_ena; // @[util.scala 28:45]
  wire  cluster_41_wea; // @[util.scala 28:45]
  wire [11:0] cluster_41_addrb; // @[util.scala 28:45]
  wire  cluster_41_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_41_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_41_doutb; // @[util.scala 28:45]
  wire  cluster_41_enb; // @[util.scala 28:45]
  wire  cluster_41_web; // @[util.scala 28:45]
  wire [11:0] cluster_42_addra; // @[util.scala 28:45]
  wire  cluster_42_clka; // @[util.scala 28:45]
  wire [47:0] cluster_42_dina; // @[util.scala 28:45]
  wire [47:0] cluster_42_douta; // @[util.scala 28:45]
  wire  cluster_42_ena; // @[util.scala 28:45]
  wire  cluster_42_wea; // @[util.scala 28:45]
  wire [11:0] cluster_42_addrb; // @[util.scala 28:45]
  wire  cluster_42_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_42_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_42_doutb; // @[util.scala 28:45]
  wire  cluster_42_enb; // @[util.scala 28:45]
  wire  cluster_42_web; // @[util.scala 28:45]
  wire [11:0] cluster_43_addra; // @[util.scala 28:45]
  wire  cluster_43_clka; // @[util.scala 28:45]
  wire [47:0] cluster_43_dina; // @[util.scala 28:45]
  wire [47:0] cluster_43_douta; // @[util.scala 28:45]
  wire  cluster_43_ena; // @[util.scala 28:45]
  wire  cluster_43_wea; // @[util.scala 28:45]
  wire [11:0] cluster_43_addrb; // @[util.scala 28:45]
  wire  cluster_43_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_43_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_43_doutb; // @[util.scala 28:45]
  wire  cluster_43_enb; // @[util.scala 28:45]
  wire  cluster_43_web; // @[util.scala 28:45]
  wire [11:0] cluster_44_addra; // @[util.scala 28:45]
  wire  cluster_44_clka; // @[util.scala 28:45]
  wire [47:0] cluster_44_dina; // @[util.scala 28:45]
  wire [47:0] cluster_44_douta; // @[util.scala 28:45]
  wire  cluster_44_ena; // @[util.scala 28:45]
  wire  cluster_44_wea; // @[util.scala 28:45]
  wire [11:0] cluster_44_addrb; // @[util.scala 28:45]
  wire  cluster_44_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_44_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_44_doutb; // @[util.scala 28:45]
  wire  cluster_44_enb; // @[util.scala 28:45]
  wire  cluster_44_web; // @[util.scala 28:45]
  wire [11:0] cluster_45_addra; // @[util.scala 28:45]
  wire  cluster_45_clka; // @[util.scala 28:45]
  wire [47:0] cluster_45_dina; // @[util.scala 28:45]
  wire [47:0] cluster_45_douta; // @[util.scala 28:45]
  wire  cluster_45_ena; // @[util.scala 28:45]
  wire  cluster_45_wea; // @[util.scala 28:45]
  wire [11:0] cluster_45_addrb; // @[util.scala 28:45]
  wire  cluster_45_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_45_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_45_doutb; // @[util.scala 28:45]
  wire  cluster_45_enb; // @[util.scala 28:45]
  wire  cluster_45_web; // @[util.scala 28:45]
  wire [11:0] cluster_46_addra; // @[util.scala 28:45]
  wire  cluster_46_clka; // @[util.scala 28:45]
  wire [47:0] cluster_46_dina; // @[util.scala 28:45]
  wire [47:0] cluster_46_douta; // @[util.scala 28:45]
  wire  cluster_46_ena; // @[util.scala 28:45]
  wire  cluster_46_wea; // @[util.scala 28:45]
  wire [11:0] cluster_46_addrb; // @[util.scala 28:45]
  wire  cluster_46_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_46_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_46_doutb; // @[util.scala 28:45]
  wire  cluster_46_enb; // @[util.scala 28:45]
  wire  cluster_46_web; // @[util.scala 28:45]
  wire [11:0] cluster_47_addra; // @[util.scala 28:45]
  wire  cluster_47_clka; // @[util.scala 28:45]
  wire [47:0] cluster_47_dina; // @[util.scala 28:45]
  wire [47:0] cluster_47_douta; // @[util.scala 28:45]
  wire  cluster_47_ena; // @[util.scala 28:45]
  wire  cluster_47_wea; // @[util.scala 28:45]
  wire [11:0] cluster_47_addrb; // @[util.scala 28:45]
  wire  cluster_47_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_47_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_47_doutb; // @[util.scala 28:45]
  wire  cluster_47_enb; // @[util.scala 28:45]
  wire  cluster_47_web; // @[util.scala 28:45]
  wire [11:0] cluster_48_addra; // @[util.scala 28:45]
  wire  cluster_48_clka; // @[util.scala 28:45]
  wire [47:0] cluster_48_dina; // @[util.scala 28:45]
  wire [47:0] cluster_48_douta; // @[util.scala 28:45]
  wire  cluster_48_ena; // @[util.scala 28:45]
  wire  cluster_48_wea; // @[util.scala 28:45]
  wire [11:0] cluster_48_addrb; // @[util.scala 28:45]
  wire  cluster_48_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_48_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_48_doutb; // @[util.scala 28:45]
  wire  cluster_48_enb; // @[util.scala 28:45]
  wire  cluster_48_web; // @[util.scala 28:45]
  wire [11:0] cluster_49_addra; // @[util.scala 28:45]
  wire  cluster_49_clka; // @[util.scala 28:45]
  wire [47:0] cluster_49_dina; // @[util.scala 28:45]
  wire [47:0] cluster_49_douta; // @[util.scala 28:45]
  wire  cluster_49_ena; // @[util.scala 28:45]
  wire  cluster_49_wea; // @[util.scala 28:45]
  wire [11:0] cluster_49_addrb; // @[util.scala 28:45]
  wire  cluster_49_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_49_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_49_doutb; // @[util.scala 28:45]
  wire  cluster_49_enb; // @[util.scala 28:45]
  wire  cluster_49_web; // @[util.scala 28:45]
  wire [11:0] cluster_50_addra; // @[util.scala 28:45]
  wire  cluster_50_clka; // @[util.scala 28:45]
  wire [47:0] cluster_50_dina; // @[util.scala 28:45]
  wire [47:0] cluster_50_douta; // @[util.scala 28:45]
  wire  cluster_50_ena; // @[util.scala 28:45]
  wire  cluster_50_wea; // @[util.scala 28:45]
  wire [11:0] cluster_50_addrb; // @[util.scala 28:45]
  wire  cluster_50_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_50_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_50_doutb; // @[util.scala 28:45]
  wire  cluster_50_enb; // @[util.scala 28:45]
  wire  cluster_50_web; // @[util.scala 28:45]
  wire [11:0] cluster_51_addra; // @[util.scala 28:45]
  wire  cluster_51_clka; // @[util.scala 28:45]
  wire [47:0] cluster_51_dina; // @[util.scala 28:45]
  wire [47:0] cluster_51_douta; // @[util.scala 28:45]
  wire  cluster_51_ena; // @[util.scala 28:45]
  wire  cluster_51_wea; // @[util.scala 28:45]
  wire [11:0] cluster_51_addrb; // @[util.scala 28:45]
  wire  cluster_51_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_51_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_51_doutb; // @[util.scala 28:45]
  wire  cluster_51_enb; // @[util.scala 28:45]
  wire  cluster_51_web; // @[util.scala 28:45]
  wire [11:0] cluster_52_addra; // @[util.scala 28:45]
  wire  cluster_52_clka; // @[util.scala 28:45]
  wire [47:0] cluster_52_dina; // @[util.scala 28:45]
  wire [47:0] cluster_52_douta; // @[util.scala 28:45]
  wire  cluster_52_ena; // @[util.scala 28:45]
  wire  cluster_52_wea; // @[util.scala 28:45]
  wire [11:0] cluster_52_addrb; // @[util.scala 28:45]
  wire  cluster_52_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_52_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_52_doutb; // @[util.scala 28:45]
  wire  cluster_52_enb; // @[util.scala 28:45]
  wire  cluster_52_web; // @[util.scala 28:45]
  wire [11:0] cluster_53_addra; // @[util.scala 28:45]
  wire  cluster_53_clka; // @[util.scala 28:45]
  wire [47:0] cluster_53_dina; // @[util.scala 28:45]
  wire [47:0] cluster_53_douta; // @[util.scala 28:45]
  wire  cluster_53_ena; // @[util.scala 28:45]
  wire  cluster_53_wea; // @[util.scala 28:45]
  wire [11:0] cluster_53_addrb; // @[util.scala 28:45]
  wire  cluster_53_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_53_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_53_doutb; // @[util.scala 28:45]
  wire  cluster_53_enb; // @[util.scala 28:45]
  wire  cluster_53_web; // @[util.scala 28:45]
  wire [11:0] cluster_54_addra; // @[util.scala 28:45]
  wire  cluster_54_clka; // @[util.scala 28:45]
  wire [47:0] cluster_54_dina; // @[util.scala 28:45]
  wire [47:0] cluster_54_douta; // @[util.scala 28:45]
  wire  cluster_54_ena; // @[util.scala 28:45]
  wire  cluster_54_wea; // @[util.scala 28:45]
  wire [11:0] cluster_54_addrb; // @[util.scala 28:45]
  wire  cluster_54_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_54_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_54_doutb; // @[util.scala 28:45]
  wire  cluster_54_enb; // @[util.scala 28:45]
  wire  cluster_54_web; // @[util.scala 28:45]
  wire [11:0] cluster_55_addra; // @[util.scala 28:45]
  wire  cluster_55_clka; // @[util.scala 28:45]
  wire [47:0] cluster_55_dina; // @[util.scala 28:45]
  wire [47:0] cluster_55_douta; // @[util.scala 28:45]
  wire  cluster_55_ena; // @[util.scala 28:45]
  wire  cluster_55_wea; // @[util.scala 28:45]
  wire [11:0] cluster_55_addrb; // @[util.scala 28:45]
  wire  cluster_55_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_55_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_55_doutb; // @[util.scala 28:45]
  wire  cluster_55_enb; // @[util.scala 28:45]
  wire  cluster_55_web; // @[util.scala 28:45]
  wire [11:0] cluster_56_addra; // @[util.scala 28:45]
  wire  cluster_56_clka; // @[util.scala 28:45]
  wire [47:0] cluster_56_dina; // @[util.scala 28:45]
  wire [47:0] cluster_56_douta; // @[util.scala 28:45]
  wire  cluster_56_ena; // @[util.scala 28:45]
  wire  cluster_56_wea; // @[util.scala 28:45]
  wire [11:0] cluster_56_addrb; // @[util.scala 28:45]
  wire  cluster_56_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_56_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_56_doutb; // @[util.scala 28:45]
  wire  cluster_56_enb; // @[util.scala 28:45]
  wire  cluster_56_web; // @[util.scala 28:45]
  wire [11:0] cluster_57_addra; // @[util.scala 28:45]
  wire  cluster_57_clka; // @[util.scala 28:45]
  wire [47:0] cluster_57_dina; // @[util.scala 28:45]
  wire [47:0] cluster_57_douta; // @[util.scala 28:45]
  wire  cluster_57_ena; // @[util.scala 28:45]
  wire  cluster_57_wea; // @[util.scala 28:45]
  wire [11:0] cluster_57_addrb; // @[util.scala 28:45]
  wire  cluster_57_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_57_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_57_doutb; // @[util.scala 28:45]
  wire  cluster_57_enb; // @[util.scala 28:45]
  wire  cluster_57_web; // @[util.scala 28:45]
  wire [11:0] cluster_58_addra; // @[util.scala 28:45]
  wire  cluster_58_clka; // @[util.scala 28:45]
  wire [47:0] cluster_58_dina; // @[util.scala 28:45]
  wire [47:0] cluster_58_douta; // @[util.scala 28:45]
  wire  cluster_58_ena; // @[util.scala 28:45]
  wire  cluster_58_wea; // @[util.scala 28:45]
  wire [11:0] cluster_58_addrb; // @[util.scala 28:45]
  wire  cluster_58_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_58_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_58_doutb; // @[util.scala 28:45]
  wire  cluster_58_enb; // @[util.scala 28:45]
  wire  cluster_58_web; // @[util.scala 28:45]
  wire [11:0] cluster_59_addra; // @[util.scala 28:45]
  wire  cluster_59_clka; // @[util.scala 28:45]
  wire [47:0] cluster_59_dina; // @[util.scala 28:45]
  wire [47:0] cluster_59_douta; // @[util.scala 28:45]
  wire  cluster_59_ena; // @[util.scala 28:45]
  wire  cluster_59_wea; // @[util.scala 28:45]
  wire [11:0] cluster_59_addrb; // @[util.scala 28:45]
  wire  cluster_59_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_59_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_59_doutb; // @[util.scala 28:45]
  wire  cluster_59_enb; // @[util.scala 28:45]
  wire  cluster_59_web; // @[util.scala 28:45]
  wire [11:0] cluster_60_addra; // @[util.scala 28:45]
  wire  cluster_60_clka; // @[util.scala 28:45]
  wire [47:0] cluster_60_dina; // @[util.scala 28:45]
  wire [47:0] cluster_60_douta; // @[util.scala 28:45]
  wire  cluster_60_ena; // @[util.scala 28:45]
  wire  cluster_60_wea; // @[util.scala 28:45]
  wire [11:0] cluster_60_addrb; // @[util.scala 28:45]
  wire  cluster_60_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_60_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_60_doutb; // @[util.scala 28:45]
  wire  cluster_60_enb; // @[util.scala 28:45]
  wire  cluster_60_web; // @[util.scala 28:45]
  wire [11:0] cluster_61_addra; // @[util.scala 28:45]
  wire  cluster_61_clka; // @[util.scala 28:45]
  wire [47:0] cluster_61_dina; // @[util.scala 28:45]
  wire [47:0] cluster_61_douta; // @[util.scala 28:45]
  wire  cluster_61_ena; // @[util.scala 28:45]
  wire  cluster_61_wea; // @[util.scala 28:45]
  wire [11:0] cluster_61_addrb; // @[util.scala 28:45]
  wire  cluster_61_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_61_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_61_doutb; // @[util.scala 28:45]
  wire  cluster_61_enb; // @[util.scala 28:45]
  wire  cluster_61_web; // @[util.scala 28:45]
  wire [11:0] cluster_62_addra; // @[util.scala 28:45]
  wire  cluster_62_clka; // @[util.scala 28:45]
  wire [47:0] cluster_62_dina; // @[util.scala 28:45]
  wire [47:0] cluster_62_douta; // @[util.scala 28:45]
  wire  cluster_62_ena; // @[util.scala 28:45]
  wire  cluster_62_wea; // @[util.scala 28:45]
  wire [11:0] cluster_62_addrb; // @[util.scala 28:45]
  wire  cluster_62_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_62_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_62_doutb; // @[util.scala 28:45]
  wire  cluster_62_enb; // @[util.scala 28:45]
  wire  cluster_62_web; // @[util.scala 28:45]
  wire [11:0] cluster_63_addra; // @[util.scala 28:45]
  wire  cluster_63_clka; // @[util.scala 28:45]
  wire [47:0] cluster_63_dina; // @[util.scala 28:45]
  wire [47:0] cluster_63_douta; // @[util.scala 28:45]
  wire  cluster_63_ena; // @[util.scala 28:45]
  wire  cluster_63_wea; // @[util.scala 28:45]
  wire [11:0] cluster_63_addrb; // @[util.scala 28:45]
  wire  cluster_63_clkb; // @[util.scala 28:45]
  wire [47:0] cluster_63_dinb; // @[util.scala 28:45]
  wire [47:0] cluster_63_doutb; // @[util.scala 28:45]
  wire  cluster_63_enb; // @[util.scala 28:45]
  wire  cluster_63_web; // @[util.scala 28:45]
  wire [17:0] _cluster_0_io_web_T = {{12'd0}, io_addrb[17:12]}; // @[util.scala 42:55]
  wire  _cluster_0_io_web_T_1 = 18'h0 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [17:0] _cluster_0_io_wea_T = {{12'd0}, io_addra[17:12]}; // @[util.scala 43:55]
  wire [47:0] doutb_0 = _cluster_0_io_web_T_1 ? cluster_0_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_1_io_web_T_1 = 18'h1 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_1 = _cluster_1_io_web_T_1 ? cluster_1_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_2_io_web_T_1 = 18'h2 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_2 = _cluster_2_io_web_T_1 ? cluster_2_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_3_io_web_T_1 = 18'h3 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_3 = _cluster_3_io_web_T_1 ? cluster_3_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_4_io_web_T_1 = 18'h4 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_4 = _cluster_4_io_web_T_1 ? cluster_4_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_5_io_web_T_1 = 18'h5 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_5 = _cluster_5_io_web_T_1 ? cluster_5_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_6_io_web_T_1 = 18'h6 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_6 = _cluster_6_io_web_T_1 ? cluster_6_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_7_io_web_T_1 = 18'h7 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_7 = _cluster_7_io_web_T_1 ? cluster_7_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_8_io_web_T_1 = 18'h8 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_8 = _cluster_8_io_web_T_1 ? cluster_8_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_9_io_web_T_1 = 18'h9 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_9 = _cluster_9_io_web_T_1 ? cluster_9_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_10_io_web_T_1 = 18'ha == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_10 = _cluster_10_io_web_T_1 ? cluster_10_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_11_io_web_T_1 = 18'hb == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_11 = _cluster_11_io_web_T_1 ? cluster_11_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_12_io_web_T_1 = 18'hc == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_12 = _cluster_12_io_web_T_1 ? cluster_12_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_13_io_web_T_1 = 18'hd == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_13 = _cluster_13_io_web_T_1 ? cluster_13_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_14_io_web_T_1 = 18'he == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_14 = _cluster_14_io_web_T_1 ? cluster_14_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_15_io_web_T_1 = 18'hf == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_15 = _cluster_15_io_web_T_1 ? cluster_15_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_16_io_web_T_1 = 18'h10 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_16 = _cluster_16_io_web_T_1 ? cluster_16_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_17_io_web_T_1 = 18'h11 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_17 = _cluster_17_io_web_T_1 ? cluster_17_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_18_io_web_T_1 = 18'h12 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_18 = _cluster_18_io_web_T_1 ? cluster_18_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_19_io_web_T_1 = 18'h13 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_19 = _cluster_19_io_web_T_1 ? cluster_19_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_20_io_web_T_1 = 18'h14 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_20 = _cluster_20_io_web_T_1 ? cluster_20_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_21_io_web_T_1 = 18'h15 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_21 = _cluster_21_io_web_T_1 ? cluster_21_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_22_io_web_T_1 = 18'h16 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_22 = _cluster_22_io_web_T_1 ? cluster_22_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_23_io_web_T_1 = 18'h17 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_23 = _cluster_23_io_web_T_1 ? cluster_23_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_24_io_web_T_1 = 18'h18 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_24 = _cluster_24_io_web_T_1 ? cluster_24_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_25_io_web_T_1 = 18'h19 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_25 = _cluster_25_io_web_T_1 ? cluster_25_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_26_io_web_T_1 = 18'h1a == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_26 = _cluster_26_io_web_T_1 ? cluster_26_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_27_io_web_T_1 = 18'h1b == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_27 = _cluster_27_io_web_T_1 ? cluster_27_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_28_io_web_T_1 = 18'h1c == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_28 = _cluster_28_io_web_T_1 ? cluster_28_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_29_io_web_T_1 = 18'h1d == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_29 = _cluster_29_io_web_T_1 ? cluster_29_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_30_io_web_T_1 = 18'h1e == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_30 = _cluster_30_io_web_T_1 ? cluster_30_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_31_io_web_T_1 = 18'h1f == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_31 = _cluster_31_io_web_T_1 ? cluster_31_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_32_io_web_T_1 = 18'h20 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_32 = _cluster_32_io_web_T_1 ? cluster_32_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_33_io_web_T_1 = 18'h21 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_33 = _cluster_33_io_web_T_1 ? cluster_33_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_34_io_web_T_1 = 18'h22 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_34 = _cluster_34_io_web_T_1 ? cluster_34_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_35_io_web_T_1 = 18'h23 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_35 = _cluster_35_io_web_T_1 ? cluster_35_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_36_io_web_T_1 = 18'h24 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_36 = _cluster_36_io_web_T_1 ? cluster_36_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_37_io_web_T_1 = 18'h25 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_37 = _cluster_37_io_web_T_1 ? cluster_37_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_38_io_web_T_1 = 18'h26 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_38 = _cluster_38_io_web_T_1 ? cluster_38_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_39_io_web_T_1 = 18'h27 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_39 = _cluster_39_io_web_T_1 ? cluster_39_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_40_io_web_T_1 = 18'h28 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_40 = _cluster_40_io_web_T_1 ? cluster_40_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_41_io_web_T_1 = 18'h29 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_41 = _cluster_41_io_web_T_1 ? cluster_41_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_42_io_web_T_1 = 18'h2a == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_42 = _cluster_42_io_web_T_1 ? cluster_42_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_43_io_web_T_1 = 18'h2b == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_43 = _cluster_43_io_web_T_1 ? cluster_43_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_44_io_web_T_1 = 18'h2c == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_44 = _cluster_44_io_web_T_1 ? cluster_44_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_45_io_web_T_1 = 18'h2d == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_45 = _cluster_45_io_web_T_1 ? cluster_45_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_46_io_web_T_1 = 18'h2e == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_46 = _cluster_46_io_web_T_1 ? cluster_46_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_47_io_web_T_1 = 18'h2f == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_47 = _cluster_47_io_web_T_1 ? cluster_47_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_48_io_web_T_1 = 18'h30 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_48 = _cluster_48_io_web_T_1 ? cluster_48_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_49_io_web_T_1 = 18'h31 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_49 = _cluster_49_io_web_T_1 ? cluster_49_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_50_io_web_T_1 = 18'h32 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_50 = _cluster_50_io_web_T_1 ? cluster_50_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_51_io_web_T_1 = 18'h33 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_51 = _cluster_51_io_web_T_1 ? cluster_51_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_52_io_web_T_1 = 18'h34 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_52 = _cluster_52_io_web_T_1 ? cluster_52_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_53_io_web_T_1 = 18'h35 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_53 = _cluster_53_io_web_T_1 ? cluster_53_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_54_io_web_T_1 = 18'h36 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_54 = _cluster_54_io_web_T_1 ? cluster_54_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_55_io_web_T_1 = 18'h37 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_55 = _cluster_55_io_web_T_1 ? cluster_55_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_56_io_web_T_1 = 18'h38 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_56 = _cluster_56_io_web_T_1 ? cluster_56_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_57_io_web_T_1 = 18'h39 == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_57 = _cluster_57_io_web_T_1 ? cluster_57_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_58_io_web_T_1 = 18'h3a == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_58 = _cluster_58_io_web_T_1 ? cluster_58_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_59_io_web_T_1 = 18'h3b == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_59 = _cluster_59_io_web_T_1 ? cluster_59_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_60_io_web_T_1 = 18'h3c == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_60 = _cluster_60_io_web_T_1 ? cluster_60_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_61_io_web_T_1 = 18'h3d == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_61 = _cluster_61_io_web_T_1 ? cluster_61_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_62_io_web_T_1 = 18'h3e == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_62 = _cluster_62_io_web_T_1 ? cluster_62_doutb : 48'h0; // @[util.scala 44:22]
  wire  _cluster_63_io_web_T_1 = 18'h3f == _cluster_0_io_web_T; // @[util.scala 42:41]
  wire [47:0] doutb_63 = _cluster_63_io_web_T_1 ? cluster_63_doutb : 48'h0; // @[util.scala 44:22]
  wire [47:0] _io_doutb_T = doutb_0 | doutb_1; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_1 = _io_doutb_T | doutb_2; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_2 = _io_doutb_T_1 | doutb_3; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_3 = _io_doutb_T_2 | doutb_4; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_4 = _io_doutb_T_3 | doutb_5; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_5 = _io_doutb_T_4 | doutb_6; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_6 = _io_doutb_T_5 | doutb_7; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_7 = _io_doutb_T_6 | doutb_8; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_8 = _io_doutb_T_7 | doutb_9; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_9 = _io_doutb_T_8 | doutb_10; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_10 = _io_doutb_T_9 | doutb_11; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_11 = _io_doutb_T_10 | doutb_12; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_12 = _io_doutb_T_11 | doutb_13; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_13 = _io_doutb_T_12 | doutb_14; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_14 = _io_doutb_T_13 | doutb_15; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_15 = _io_doutb_T_14 | doutb_16; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_16 = _io_doutb_T_15 | doutb_17; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_17 = _io_doutb_T_16 | doutb_18; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_18 = _io_doutb_T_17 | doutb_19; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_19 = _io_doutb_T_18 | doutb_20; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_20 = _io_doutb_T_19 | doutb_21; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_21 = _io_doutb_T_20 | doutb_22; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_22 = _io_doutb_T_21 | doutb_23; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_23 = _io_doutb_T_22 | doutb_24; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_24 = _io_doutb_T_23 | doutb_25; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_25 = _io_doutb_T_24 | doutb_26; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_26 = _io_doutb_T_25 | doutb_27; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_27 = _io_doutb_T_26 | doutb_28; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_28 = _io_doutb_T_27 | doutb_29; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_29 = _io_doutb_T_28 | doutb_30; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_30 = _io_doutb_T_29 | doutb_31; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_31 = _io_doutb_T_30 | doutb_32; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_32 = _io_doutb_T_31 | doutb_33; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_33 = _io_doutb_T_32 | doutb_34; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_34 = _io_doutb_T_33 | doutb_35; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_35 = _io_doutb_T_34 | doutb_36; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_36 = _io_doutb_T_35 | doutb_37; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_37 = _io_doutb_T_36 | doutb_38; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_38 = _io_doutb_T_37 | doutb_39; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_39 = _io_doutb_T_38 | doutb_40; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_40 = _io_doutb_T_39 | doutb_41; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_41 = _io_doutb_T_40 | doutb_42; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_42 = _io_doutb_T_41 | doutb_43; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_43 = _io_doutb_T_42 | doutb_44; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_44 = _io_doutb_T_43 | doutb_45; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_45 = _io_doutb_T_44 | doutb_46; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_46 = _io_doutb_T_45 | doutb_47; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_47 = _io_doutb_T_46 | doutb_48; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_48 = _io_doutb_T_47 | doutb_49; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_49 = _io_doutb_T_48 | doutb_50; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_50 = _io_doutb_T_49 | doutb_51; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_51 = _io_doutb_T_50 | doutb_52; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_52 = _io_doutb_T_51 | doutb_53; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_53 = _io_doutb_T_52 | doutb_54; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_54 = _io_doutb_T_53 | doutb_55; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_55 = _io_doutb_T_54 | doutb_56; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_56 = _io_doutb_T_55 | doutb_57; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_57 = _io_doutb_T_56 | doutb_58; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_58 = _io_doutb_T_57 | doutb_59; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_59 = _io_doutb_T_58 | doutb_60; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_60 = _io_doutb_T_59 | doutb_61; // @[util.scala 49:29]
  wire [47:0] _io_doutb_T_61 = _io_doutb_T_60 | doutb_62; // @[util.scala 49:29]
  URAM cluster_0 ( // @[util.scala 28:45]
    .addra(cluster_0_addra),
    .clka(cluster_0_clka),
    .dina(cluster_0_dina),
    .douta(cluster_0_douta),
    .ena(cluster_0_ena),
    .wea(cluster_0_wea),
    .addrb(cluster_0_addrb),
    .clkb(cluster_0_clkb),
    .dinb(cluster_0_dinb),
    .doutb(cluster_0_doutb),
    .enb(cluster_0_enb),
    .web(cluster_0_web)
  );
  URAM cluster_1 ( // @[util.scala 28:45]
    .addra(cluster_1_addra),
    .clka(cluster_1_clka),
    .dina(cluster_1_dina),
    .douta(cluster_1_douta),
    .ena(cluster_1_ena),
    .wea(cluster_1_wea),
    .addrb(cluster_1_addrb),
    .clkb(cluster_1_clkb),
    .dinb(cluster_1_dinb),
    .doutb(cluster_1_doutb),
    .enb(cluster_1_enb),
    .web(cluster_1_web)
  );
  URAM cluster_2 ( // @[util.scala 28:45]
    .addra(cluster_2_addra),
    .clka(cluster_2_clka),
    .dina(cluster_2_dina),
    .douta(cluster_2_douta),
    .ena(cluster_2_ena),
    .wea(cluster_2_wea),
    .addrb(cluster_2_addrb),
    .clkb(cluster_2_clkb),
    .dinb(cluster_2_dinb),
    .doutb(cluster_2_doutb),
    .enb(cluster_2_enb),
    .web(cluster_2_web)
  );
  URAM cluster_3 ( // @[util.scala 28:45]
    .addra(cluster_3_addra),
    .clka(cluster_3_clka),
    .dina(cluster_3_dina),
    .douta(cluster_3_douta),
    .ena(cluster_3_ena),
    .wea(cluster_3_wea),
    .addrb(cluster_3_addrb),
    .clkb(cluster_3_clkb),
    .dinb(cluster_3_dinb),
    .doutb(cluster_3_doutb),
    .enb(cluster_3_enb),
    .web(cluster_3_web)
  );
  URAM cluster_4 ( // @[util.scala 28:45]
    .addra(cluster_4_addra),
    .clka(cluster_4_clka),
    .dina(cluster_4_dina),
    .douta(cluster_4_douta),
    .ena(cluster_4_ena),
    .wea(cluster_4_wea),
    .addrb(cluster_4_addrb),
    .clkb(cluster_4_clkb),
    .dinb(cluster_4_dinb),
    .doutb(cluster_4_doutb),
    .enb(cluster_4_enb),
    .web(cluster_4_web)
  );
  URAM cluster_5 ( // @[util.scala 28:45]
    .addra(cluster_5_addra),
    .clka(cluster_5_clka),
    .dina(cluster_5_dina),
    .douta(cluster_5_douta),
    .ena(cluster_5_ena),
    .wea(cluster_5_wea),
    .addrb(cluster_5_addrb),
    .clkb(cluster_5_clkb),
    .dinb(cluster_5_dinb),
    .doutb(cluster_5_doutb),
    .enb(cluster_5_enb),
    .web(cluster_5_web)
  );
  URAM cluster_6 ( // @[util.scala 28:45]
    .addra(cluster_6_addra),
    .clka(cluster_6_clka),
    .dina(cluster_6_dina),
    .douta(cluster_6_douta),
    .ena(cluster_6_ena),
    .wea(cluster_6_wea),
    .addrb(cluster_6_addrb),
    .clkb(cluster_6_clkb),
    .dinb(cluster_6_dinb),
    .doutb(cluster_6_doutb),
    .enb(cluster_6_enb),
    .web(cluster_6_web)
  );
  URAM cluster_7 ( // @[util.scala 28:45]
    .addra(cluster_7_addra),
    .clka(cluster_7_clka),
    .dina(cluster_7_dina),
    .douta(cluster_7_douta),
    .ena(cluster_7_ena),
    .wea(cluster_7_wea),
    .addrb(cluster_7_addrb),
    .clkb(cluster_7_clkb),
    .dinb(cluster_7_dinb),
    .doutb(cluster_7_doutb),
    .enb(cluster_7_enb),
    .web(cluster_7_web)
  );
  URAM cluster_8 ( // @[util.scala 28:45]
    .addra(cluster_8_addra),
    .clka(cluster_8_clka),
    .dina(cluster_8_dina),
    .douta(cluster_8_douta),
    .ena(cluster_8_ena),
    .wea(cluster_8_wea),
    .addrb(cluster_8_addrb),
    .clkb(cluster_8_clkb),
    .dinb(cluster_8_dinb),
    .doutb(cluster_8_doutb),
    .enb(cluster_8_enb),
    .web(cluster_8_web)
  );
  URAM cluster_9 ( // @[util.scala 28:45]
    .addra(cluster_9_addra),
    .clka(cluster_9_clka),
    .dina(cluster_9_dina),
    .douta(cluster_9_douta),
    .ena(cluster_9_ena),
    .wea(cluster_9_wea),
    .addrb(cluster_9_addrb),
    .clkb(cluster_9_clkb),
    .dinb(cluster_9_dinb),
    .doutb(cluster_9_doutb),
    .enb(cluster_9_enb),
    .web(cluster_9_web)
  );
  URAM cluster_10 ( // @[util.scala 28:45]
    .addra(cluster_10_addra),
    .clka(cluster_10_clka),
    .dina(cluster_10_dina),
    .douta(cluster_10_douta),
    .ena(cluster_10_ena),
    .wea(cluster_10_wea),
    .addrb(cluster_10_addrb),
    .clkb(cluster_10_clkb),
    .dinb(cluster_10_dinb),
    .doutb(cluster_10_doutb),
    .enb(cluster_10_enb),
    .web(cluster_10_web)
  );
  URAM cluster_11 ( // @[util.scala 28:45]
    .addra(cluster_11_addra),
    .clka(cluster_11_clka),
    .dina(cluster_11_dina),
    .douta(cluster_11_douta),
    .ena(cluster_11_ena),
    .wea(cluster_11_wea),
    .addrb(cluster_11_addrb),
    .clkb(cluster_11_clkb),
    .dinb(cluster_11_dinb),
    .doutb(cluster_11_doutb),
    .enb(cluster_11_enb),
    .web(cluster_11_web)
  );
  URAM cluster_12 ( // @[util.scala 28:45]
    .addra(cluster_12_addra),
    .clka(cluster_12_clka),
    .dina(cluster_12_dina),
    .douta(cluster_12_douta),
    .ena(cluster_12_ena),
    .wea(cluster_12_wea),
    .addrb(cluster_12_addrb),
    .clkb(cluster_12_clkb),
    .dinb(cluster_12_dinb),
    .doutb(cluster_12_doutb),
    .enb(cluster_12_enb),
    .web(cluster_12_web)
  );
  URAM cluster_13 ( // @[util.scala 28:45]
    .addra(cluster_13_addra),
    .clka(cluster_13_clka),
    .dina(cluster_13_dina),
    .douta(cluster_13_douta),
    .ena(cluster_13_ena),
    .wea(cluster_13_wea),
    .addrb(cluster_13_addrb),
    .clkb(cluster_13_clkb),
    .dinb(cluster_13_dinb),
    .doutb(cluster_13_doutb),
    .enb(cluster_13_enb),
    .web(cluster_13_web)
  );
  URAM cluster_14 ( // @[util.scala 28:45]
    .addra(cluster_14_addra),
    .clka(cluster_14_clka),
    .dina(cluster_14_dina),
    .douta(cluster_14_douta),
    .ena(cluster_14_ena),
    .wea(cluster_14_wea),
    .addrb(cluster_14_addrb),
    .clkb(cluster_14_clkb),
    .dinb(cluster_14_dinb),
    .doutb(cluster_14_doutb),
    .enb(cluster_14_enb),
    .web(cluster_14_web)
  );
  URAM cluster_15 ( // @[util.scala 28:45]
    .addra(cluster_15_addra),
    .clka(cluster_15_clka),
    .dina(cluster_15_dina),
    .douta(cluster_15_douta),
    .ena(cluster_15_ena),
    .wea(cluster_15_wea),
    .addrb(cluster_15_addrb),
    .clkb(cluster_15_clkb),
    .dinb(cluster_15_dinb),
    .doutb(cluster_15_doutb),
    .enb(cluster_15_enb),
    .web(cluster_15_web)
  );
  URAM cluster_16 ( // @[util.scala 28:45]
    .addra(cluster_16_addra),
    .clka(cluster_16_clka),
    .dina(cluster_16_dina),
    .douta(cluster_16_douta),
    .ena(cluster_16_ena),
    .wea(cluster_16_wea),
    .addrb(cluster_16_addrb),
    .clkb(cluster_16_clkb),
    .dinb(cluster_16_dinb),
    .doutb(cluster_16_doutb),
    .enb(cluster_16_enb),
    .web(cluster_16_web)
  );
  URAM cluster_17 ( // @[util.scala 28:45]
    .addra(cluster_17_addra),
    .clka(cluster_17_clka),
    .dina(cluster_17_dina),
    .douta(cluster_17_douta),
    .ena(cluster_17_ena),
    .wea(cluster_17_wea),
    .addrb(cluster_17_addrb),
    .clkb(cluster_17_clkb),
    .dinb(cluster_17_dinb),
    .doutb(cluster_17_doutb),
    .enb(cluster_17_enb),
    .web(cluster_17_web)
  );
  URAM cluster_18 ( // @[util.scala 28:45]
    .addra(cluster_18_addra),
    .clka(cluster_18_clka),
    .dina(cluster_18_dina),
    .douta(cluster_18_douta),
    .ena(cluster_18_ena),
    .wea(cluster_18_wea),
    .addrb(cluster_18_addrb),
    .clkb(cluster_18_clkb),
    .dinb(cluster_18_dinb),
    .doutb(cluster_18_doutb),
    .enb(cluster_18_enb),
    .web(cluster_18_web)
  );
  URAM cluster_19 ( // @[util.scala 28:45]
    .addra(cluster_19_addra),
    .clka(cluster_19_clka),
    .dina(cluster_19_dina),
    .douta(cluster_19_douta),
    .ena(cluster_19_ena),
    .wea(cluster_19_wea),
    .addrb(cluster_19_addrb),
    .clkb(cluster_19_clkb),
    .dinb(cluster_19_dinb),
    .doutb(cluster_19_doutb),
    .enb(cluster_19_enb),
    .web(cluster_19_web)
  );
  URAM cluster_20 ( // @[util.scala 28:45]
    .addra(cluster_20_addra),
    .clka(cluster_20_clka),
    .dina(cluster_20_dina),
    .douta(cluster_20_douta),
    .ena(cluster_20_ena),
    .wea(cluster_20_wea),
    .addrb(cluster_20_addrb),
    .clkb(cluster_20_clkb),
    .dinb(cluster_20_dinb),
    .doutb(cluster_20_doutb),
    .enb(cluster_20_enb),
    .web(cluster_20_web)
  );
  URAM cluster_21 ( // @[util.scala 28:45]
    .addra(cluster_21_addra),
    .clka(cluster_21_clka),
    .dina(cluster_21_dina),
    .douta(cluster_21_douta),
    .ena(cluster_21_ena),
    .wea(cluster_21_wea),
    .addrb(cluster_21_addrb),
    .clkb(cluster_21_clkb),
    .dinb(cluster_21_dinb),
    .doutb(cluster_21_doutb),
    .enb(cluster_21_enb),
    .web(cluster_21_web)
  );
  URAM cluster_22 ( // @[util.scala 28:45]
    .addra(cluster_22_addra),
    .clka(cluster_22_clka),
    .dina(cluster_22_dina),
    .douta(cluster_22_douta),
    .ena(cluster_22_ena),
    .wea(cluster_22_wea),
    .addrb(cluster_22_addrb),
    .clkb(cluster_22_clkb),
    .dinb(cluster_22_dinb),
    .doutb(cluster_22_doutb),
    .enb(cluster_22_enb),
    .web(cluster_22_web)
  );
  URAM cluster_23 ( // @[util.scala 28:45]
    .addra(cluster_23_addra),
    .clka(cluster_23_clka),
    .dina(cluster_23_dina),
    .douta(cluster_23_douta),
    .ena(cluster_23_ena),
    .wea(cluster_23_wea),
    .addrb(cluster_23_addrb),
    .clkb(cluster_23_clkb),
    .dinb(cluster_23_dinb),
    .doutb(cluster_23_doutb),
    .enb(cluster_23_enb),
    .web(cluster_23_web)
  );
  URAM cluster_24 ( // @[util.scala 28:45]
    .addra(cluster_24_addra),
    .clka(cluster_24_clka),
    .dina(cluster_24_dina),
    .douta(cluster_24_douta),
    .ena(cluster_24_ena),
    .wea(cluster_24_wea),
    .addrb(cluster_24_addrb),
    .clkb(cluster_24_clkb),
    .dinb(cluster_24_dinb),
    .doutb(cluster_24_doutb),
    .enb(cluster_24_enb),
    .web(cluster_24_web)
  );
  URAM cluster_25 ( // @[util.scala 28:45]
    .addra(cluster_25_addra),
    .clka(cluster_25_clka),
    .dina(cluster_25_dina),
    .douta(cluster_25_douta),
    .ena(cluster_25_ena),
    .wea(cluster_25_wea),
    .addrb(cluster_25_addrb),
    .clkb(cluster_25_clkb),
    .dinb(cluster_25_dinb),
    .doutb(cluster_25_doutb),
    .enb(cluster_25_enb),
    .web(cluster_25_web)
  );
  URAM cluster_26 ( // @[util.scala 28:45]
    .addra(cluster_26_addra),
    .clka(cluster_26_clka),
    .dina(cluster_26_dina),
    .douta(cluster_26_douta),
    .ena(cluster_26_ena),
    .wea(cluster_26_wea),
    .addrb(cluster_26_addrb),
    .clkb(cluster_26_clkb),
    .dinb(cluster_26_dinb),
    .doutb(cluster_26_doutb),
    .enb(cluster_26_enb),
    .web(cluster_26_web)
  );
  URAM cluster_27 ( // @[util.scala 28:45]
    .addra(cluster_27_addra),
    .clka(cluster_27_clka),
    .dina(cluster_27_dina),
    .douta(cluster_27_douta),
    .ena(cluster_27_ena),
    .wea(cluster_27_wea),
    .addrb(cluster_27_addrb),
    .clkb(cluster_27_clkb),
    .dinb(cluster_27_dinb),
    .doutb(cluster_27_doutb),
    .enb(cluster_27_enb),
    .web(cluster_27_web)
  );
  URAM cluster_28 ( // @[util.scala 28:45]
    .addra(cluster_28_addra),
    .clka(cluster_28_clka),
    .dina(cluster_28_dina),
    .douta(cluster_28_douta),
    .ena(cluster_28_ena),
    .wea(cluster_28_wea),
    .addrb(cluster_28_addrb),
    .clkb(cluster_28_clkb),
    .dinb(cluster_28_dinb),
    .doutb(cluster_28_doutb),
    .enb(cluster_28_enb),
    .web(cluster_28_web)
  );
  URAM cluster_29 ( // @[util.scala 28:45]
    .addra(cluster_29_addra),
    .clka(cluster_29_clka),
    .dina(cluster_29_dina),
    .douta(cluster_29_douta),
    .ena(cluster_29_ena),
    .wea(cluster_29_wea),
    .addrb(cluster_29_addrb),
    .clkb(cluster_29_clkb),
    .dinb(cluster_29_dinb),
    .doutb(cluster_29_doutb),
    .enb(cluster_29_enb),
    .web(cluster_29_web)
  );
  URAM cluster_30 ( // @[util.scala 28:45]
    .addra(cluster_30_addra),
    .clka(cluster_30_clka),
    .dina(cluster_30_dina),
    .douta(cluster_30_douta),
    .ena(cluster_30_ena),
    .wea(cluster_30_wea),
    .addrb(cluster_30_addrb),
    .clkb(cluster_30_clkb),
    .dinb(cluster_30_dinb),
    .doutb(cluster_30_doutb),
    .enb(cluster_30_enb),
    .web(cluster_30_web)
  );
  URAM cluster_31 ( // @[util.scala 28:45]
    .addra(cluster_31_addra),
    .clka(cluster_31_clka),
    .dina(cluster_31_dina),
    .douta(cluster_31_douta),
    .ena(cluster_31_ena),
    .wea(cluster_31_wea),
    .addrb(cluster_31_addrb),
    .clkb(cluster_31_clkb),
    .dinb(cluster_31_dinb),
    .doutb(cluster_31_doutb),
    .enb(cluster_31_enb),
    .web(cluster_31_web)
  );
  URAM cluster_32 ( // @[util.scala 28:45]
    .addra(cluster_32_addra),
    .clka(cluster_32_clka),
    .dina(cluster_32_dina),
    .douta(cluster_32_douta),
    .ena(cluster_32_ena),
    .wea(cluster_32_wea),
    .addrb(cluster_32_addrb),
    .clkb(cluster_32_clkb),
    .dinb(cluster_32_dinb),
    .doutb(cluster_32_doutb),
    .enb(cluster_32_enb),
    .web(cluster_32_web)
  );
  URAM cluster_33 ( // @[util.scala 28:45]
    .addra(cluster_33_addra),
    .clka(cluster_33_clka),
    .dina(cluster_33_dina),
    .douta(cluster_33_douta),
    .ena(cluster_33_ena),
    .wea(cluster_33_wea),
    .addrb(cluster_33_addrb),
    .clkb(cluster_33_clkb),
    .dinb(cluster_33_dinb),
    .doutb(cluster_33_doutb),
    .enb(cluster_33_enb),
    .web(cluster_33_web)
  );
  URAM cluster_34 ( // @[util.scala 28:45]
    .addra(cluster_34_addra),
    .clka(cluster_34_clka),
    .dina(cluster_34_dina),
    .douta(cluster_34_douta),
    .ena(cluster_34_ena),
    .wea(cluster_34_wea),
    .addrb(cluster_34_addrb),
    .clkb(cluster_34_clkb),
    .dinb(cluster_34_dinb),
    .doutb(cluster_34_doutb),
    .enb(cluster_34_enb),
    .web(cluster_34_web)
  );
  URAM cluster_35 ( // @[util.scala 28:45]
    .addra(cluster_35_addra),
    .clka(cluster_35_clka),
    .dina(cluster_35_dina),
    .douta(cluster_35_douta),
    .ena(cluster_35_ena),
    .wea(cluster_35_wea),
    .addrb(cluster_35_addrb),
    .clkb(cluster_35_clkb),
    .dinb(cluster_35_dinb),
    .doutb(cluster_35_doutb),
    .enb(cluster_35_enb),
    .web(cluster_35_web)
  );
  URAM cluster_36 ( // @[util.scala 28:45]
    .addra(cluster_36_addra),
    .clka(cluster_36_clka),
    .dina(cluster_36_dina),
    .douta(cluster_36_douta),
    .ena(cluster_36_ena),
    .wea(cluster_36_wea),
    .addrb(cluster_36_addrb),
    .clkb(cluster_36_clkb),
    .dinb(cluster_36_dinb),
    .doutb(cluster_36_doutb),
    .enb(cluster_36_enb),
    .web(cluster_36_web)
  );
  URAM cluster_37 ( // @[util.scala 28:45]
    .addra(cluster_37_addra),
    .clka(cluster_37_clka),
    .dina(cluster_37_dina),
    .douta(cluster_37_douta),
    .ena(cluster_37_ena),
    .wea(cluster_37_wea),
    .addrb(cluster_37_addrb),
    .clkb(cluster_37_clkb),
    .dinb(cluster_37_dinb),
    .doutb(cluster_37_doutb),
    .enb(cluster_37_enb),
    .web(cluster_37_web)
  );
  URAM cluster_38 ( // @[util.scala 28:45]
    .addra(cluster_38_addra),
    .clka(cluster_38_clka),
    .dina(cluster_38_dina),
    .douta(cluster_38_douta),
    .ena(cluster_38_ena),
    .wea(cluster_38_wea),
    .addrb(cluster_38_addrb),
    .clkb(cluster_38_clkb),
    .dinb(cluster_38_dinb),
    .doutb(cluster_38_doutb),
    .enb(cluster_38_enb),
    .web(cluster_38_web)
  );
  URAM cluster_39 ( // @[util.scala 28:45]
    .addra(cluster_39_addra),
    .clka(cluster_39_clka),
    .dina(cluster_39_dina),
    .douta(cluster_39_douta),
    .ena(cluster_39_ena),
    .wea(cluster_39_wea),
    .addrb(cluster_39_addrb),
    .clkb(cluster_39_clkb),
    .dinb(cluster_39_dinb),
    .doutb(cluster_39_doutb),
    .enb(cluster_39_enb),
    .web(cluster_39_web)
  );
  URAM cluster_40 ( // @[util.scala 28:45]
    .addra(cluster_40_addra),
    .clka(cluster_40_clka),
    .dina(cluster_40_dina),
    .douta(cluster_40_douta),
    .ena(cluster_40_ena),
    .wea(cluster_40_wea),
    .addrb(cluster_40_addrb),
    .clkb(cluster_40_clkb),
    .dinb(cluster_40_dinb),
    .doutb(cluster_40_doutb),
    .enb(cluster_40_enb),
    .web(cluster_40_web)
  );
  URAM cluster_41 ( // @[util.scala 28:45]
    .addra(cluster_41_addra),
    .clka(cluster_41_clka),
    .dina(cluster_41_dina),
    .douta(cluster_41_douta),
    .ena(cluster_41_ena),
    .wea(cluster_41_wea),
    .addrb(cluster_41_addrb),
    .clkb(cluster_41_clkb),
    .dinb(cluster_41_dinb),
    .doutb(cluster_41_doutb),
    .enb(cluster_41_enb),
    .web(cluster_41_web)
  );
  URAM cluster_42 ( // @[util.scala 28:45]
    .addra(cluster_42_addra),
    .clka(cluster_42_clka),
    .dina(cluster_42_dina),
    .douta(cluster_42_douta),
    .ena(cluster_42_ena),
    .wea(cluster_42_wea),
    .addrb(cluster_42_addrb),
    .clkb(cluster_42_clkb),
    .dinb(cluster_42_dinb),
    .doutb(cluster_42_doutb),
    .enb(cluster_42_enb),
    .web(cluster_42_web)
  );
  URAM cluster_43 ( // @[util.scala 28:45]
    .addra(cluster_43_addra),
    .clka(cluster_43_clka),
    .dina(cluster_43_dina),
    .douta(cluster_43_douta),
    .ena(cluster_43_ena),
    .wea(cluster_43_wea),
    .addrb(cluster_43_addrb),
    .clkb(cluster_43_clkb),
    .dinb(cluster_43_dinb),
    .doutb(cluster_43_doutb),
    .enb(cluster_43_enb),
    .web(cluster_43_web)
  );
  URAM cluster_44 ( // @[util.scala 28:45]
    .addra(cluster_44_addra),
    .clka(cluster_44_clka),
    .dina(cluster_44_dina),
    .douta(cluster_44_douta),
    .ena(cluster_44_ena),
    .wea(cluster_44_wea),
    .addrb(cluster_44_addrb),
    .clkb(cluster_44_clkb),
    .dinb(cluster_44_dinb),
    .doutb(cluster_44_doutb),
    .enb(cluster_44_enb),
    .web(cluster_44_web)
  );
  URAM cluster_45 ( // @[util.scala 28:45]
    .addra(cluster_45_addra),
    .clka(cluster_45_clka),
    .dina(cluster_45_dina),
    .douta(cluster_45_douta),
    .ena(cluster_45_ena),
    .wea(cluster_45_wea),
    .addrb(cluster_45_addrb),
    .clkb(cluster_45_clkb),
    .dinb(cluster_45_dinb),
    .doutb(cluster_45_doutb),
    .enb(cluster_45_enb),
    .web(cluster_45_web)
  );
  URAM cluster_46 ( // @[util.scala 28:45]
    .addra(cluster_46_addra),
    .clka(cluster_46_clka),
    .dina(cluster_46_dina),
    .douta(cluster_46_douta),
    .ena(cluster_46_ena),
    .wea(cluster_46_wea),
    .addrb(cluster_46_addrb),
    .clkb(cluster_46_clkb),
    .dinb(cluster_46_dinb),
    .doutb(cluster_46_doutb),
    .enb(cluster_46_enb),
    .web(cluster_46_web)
  );
  URAM cluster_47 ( // @[util.scala 28:45]
    .addra(cluster_47_addra),
    .clka(cluster_47_clka),
    .dina(cluster_47_dina),
    .douta(cluster_47_douta),
    .ena(cluster_47_ena),
    .wea(cluster_47_wea),
    .addrb(cluster_47_addrb),
    .clkb(cluster_47_clkb),
    .dinb(cluster_47_dinb),
    .doutb(cluster_47_doutb),
    .enb(cluster_47_enb),
    .web(cluster_47_web)
  );
  URAM cluster_48 ( // @[util.scala 28:45]
    .addra(cluster_48_addra),
    .clka(cluster_48_clka),
    .dina(cluster_48_dina),
    .douta(cluster_48_douta),
    .ena(cluster_48_ena),
    .wea(cluster_48_wea),
    .addrb(cluster_48_addrb),
    .clkb(cluster_48_clkb),
    .dinb(cluster_48_dinb),
    .doutb(cluster_48_doutb),
    .enb(cluster_48_enb),
    .web(cluster_48_web)
  );
  URAM cluster_49 ( // @[util.scala 28:45]
    .addra(cluster_49_addra),
    .clka(cluster_49_clka),
    .dina(cluster_49_dina),
    .douta(cluster_49_douta),
    .ena(cluster_49_ena),
    .wea(cluster_49_wea),
    .addrb(cluster_49_addrb),
    .clkb(cluster_49_clkb),
    .dinb(cluster_49_dinb),
    .doutb(cluster_49_doutb),
    .enb(cluster_49_enb),
    .web(cluster_49_web)
  );
  URAM cluster_50 ( // @[util.scala 28:45]
    .addra(cluster_50_addra),
    .clka(cluster_50_clka),
    .dina(cluster_50_dina),
    .douta(cluster_50_douta),
    .ena(cluster_50_ena),
    .wea(cluster_50_wea),
    .addrb(cluster_50_addrb),
    .clkb(cluster_50_clkb),
    .dinb(cluster_50_dinb),
    .doutb(cluster_50_doutb),
    .enb(cluster_50_enb),
    .web(cluster_50_web)
  );
  URAM cluster_51 ( // @[util.scala 28:45]
    .addra(cluster_51_addra),
    .clka(cluster_51_clka),
    .dina(cluster_51_dina),
    .douta(cluster_51_douta),
    .ena(cluster_51_ena),
    .wea(cluster_51_wea),
    .addrb(cluster_51_addrb),
    .clkb(cluster_51_clkb),
    .dinb(cluster_51_dinb),
    .doutb(cluster_51_doutb),
    .enb(cluster_51_enb),
    .web(cluster_51_web)
  );
  URAM cluster_52 ( // @[util.scala 28:45]
    .addra(cluster_52_addra),
    .clka(cluster_52_clka),
    .dina(cluster_52_dina),
    .douta(cluster_52_douta),
    .ena(cluster_52_ena),
    .wea(cluster_52_wea),
    .addrb(cluster_52_addrb),
    .clkb(cluster_52_clkb),
    .dinb(cluster_52_dinb),
    .doutb(cluster_52_doutb),
    .enb(cluster_52_enb),
    .web(cluster_52_web)
  );
  URAM cluster_53 ( // @[util.scala 28:45]
    .addra(cluster_53_addra),
    .clka(cluster_53_clka),
    .dina(cluster_53_dina),
    .douta(cluster_53_douta),
    .ena(cluster_53_ena),
    .wea(cluster_53_wea),
    .addrb(cluster_53_addrb),
    .clkb(cluster_53_clkb),
    .dinb(cluster_53_dinb),
    .doutb(cluster_53_doutb),
    .enb(cluster_53_enb),
    .web(cluster_53_web)
  );
  URAM cluster_54 ( // @[util.scala 28:45]
    .addra(cluster_54_addra),
    .clka(cluster_54_clka),
    .dina(cluster_54_dina),
    .douta(cluster_54_douta),
    .ena(cluster_54_ena),
    .wea(cluster_54_wea),
    .addrb(cluster_54_addrb),
    .clkb(cluster_54_clkb),
    .dinb(cluster_54_dinb),
    .doutb(cluster_54_doutb),
    .enb(cluster_54_enb),
    .web(cluster_54_web)
  );
  URAM cluster_55 ( // @[util.scala 28:45]
    .addra(cluster_55_addra),
    .clka(cluster_55_clka),
    .dina(cluster_55_dina),
    .douta(cluster_55_douta),
    .ena(cluster_55_ena),
    .wea(cluster_55_wea),
    .addrb(cluster_55_addrb),
    .clkb(cluster_55_clkb),
    .dinb(cluster_55_dinb),
    .doutb(cluster_55_doutb),
    .enb(cluster_55_enb),
    .web(cluster_55_web)
  );
  URAM cluster_56 ( // @[util.scala 28:45]
    .addra(cluster_56_addra),
    .clka(cluster_56_clka),
    .dina(cluster_56_dina),
    .douta(cluster_56_douta),
    .ena(cluster_56_ena),
    .wea(cluster_56_wea),
    .addrb(cluster_56_addrb),
    .clkb(cluster_56_clkb),
    .dinb(cluster_56_dinb),
    .doutb(cluster_56_doutb),
    .enb(cluster_56_enb),
    .web(cluster_56_web)
  );
  URAM cluster_57 ( // @[util.scala 28:45]
    .addra(cluster_57_addra),
    .clka(cluster_57_clka),
    .dina(cluster_57_dina),
    .douta(cluster_57_douta),
    .ena(cluster_57_ena),
    .wea(cluster_57_wea),
    .addrb(cluster_57_addrb),
    .clkb(cluster_57_clkb),
    .dinb(cluster_57_dinb),
    .doutb(cluster_57_doutb),
    .enb(cluster_57_enb),
    .web(cluster_57_web)
  );
  URAM cluster_58 ( // @[util.scala 28:45]
    .addra(cluster_58_addra),
    .clka(cluster_58_clka),
    .dina(cluster_58_dina),
    .douta(cluster_58_douta),
    .ena(cluster_58_ena),
    .wea(cluster_58_wea),
    .addrb(cluster_58_addrb),
    .clkb(cluster_58_clkb),
    .dinb(cluster_58_dinb),
    .doutb(cluster_58_doutb),
    .enb(cluster_58_enb),
    .web(cluster_58_web)
  );
  URAM cluster_59 ( // @[util.scala 28:45]
    .addra(cluster_59_addra),
    .clka(cluster_59_clka),
    .dina(cluster_59_dina),
    .douta(cluster_59_douta),
    .ena(cluster_59_ena),
    .wea(cluster_59_wea),
    .addrb(cluster_59_addrb),
    .clkb(cluster_59_clkb),
    .dinb(cluster_59_dinb),
    .doutb(cluster_59_doutb),
    .enb(cluster_59_enb),
    .web(cluster_59_web)
  );
  URAM cluster_60 ( // @[util.scala 28:45]
    .addra(cluster_60_addra),
    .clka(cluster_60_clka),
    .dina(cluster_60_dina),
    .douta(cluster_60_douta),
    .ena(cluster_60_ena),
    .wea(cluster_60_wea),
    .addrb(cluster_60_addrb),
    .clkb(cluster_60_clkb),
    .dinb(cluster_60_dinb),
    .doutb(cluster_60_doutb),
    .enb(cluster_60_enb),
    .web(cluster_60_web)
  );
  URAM cluster_61 ( // @[util.scala 28:45]
    .addra(cluster_61_addra),
    .clka(cluster_61_clka),
    .dina(cluster_61_dina),
    .douta(cluster_61_douta),
    .ena(cluster_61_ena),
    .wea(cluster_61_wea),
    .addrb(cluster_61_addrb),
    .clkb(cluster_61_clkb),
    .dinb(cluster_61_dinb),
    .doutb(cluster_61_doutb),
    .enb(cluster_61_enb),
    .web(cluster_61_web)
  );
  URAM cluster_62 ( // @[util.scala 28:45]
    .addra(cluster_62_addra),
    .clka(cluster_62_clka),
    .dina(cluster_62_dina),
    .douta(cluster_62_douta),
    .ena(cluster_62_ena),
    .wea(cluster_62_wea),
    .addrb(cluster_62_addrb),
    .clkb(cluster_62_clkb),
    .dinb(cluster_62_dinb),
    .doutb(cluster_62_doutb),
    .enb(cluster_62_enb),
    .web(cluster_62_web)
  );
  URAM cluster_63 ( // @[util.scala 28:45]
    .addra(cluster_63_addra),
    .clka(cluster_63_clka),
    .dina(cluster_63_dina),
    .douta(cluster_63_douta),
    .ena(cluster_63_ena),
    .wea(cluster_63_wea),
    .addrb(cluster_63_addrb),
    .clkb(cluster_63_clkb),
    .dinb(cluster_63_dinb),
    .doutb(cluster_63_doutb),
    .enb(cluster_63_enb),
    .web(cluster_63_web)
  );
  assign io_doutb = _io_doutb_T_61 | doutb_63; // @[util.scala 49:29]
  assign cluster_0_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_0_clka = io_clka; // @[util.scala 35:17]
  assign cluster_0_dina = io_dina; // @[util.scala 39:17]
  assign cluster_0_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_0_wea = io_wea & 18'h0 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_0_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_0_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_0_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_0_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_0_web = 1'h0; // @[util.scala 42:26]
  assign cluster_1_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_1_clka = io_clka; // @[util.scala 35:17]
  assign cluster_1_dina = io_dina; // @[util.scala 39:17]
  assign cluster_1_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_1_wea = io_wea & 18'h1 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_1_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_1_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_1_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_1_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_1_web = 1'h0; // @[util.scala 42:26]
  assign cluster_2_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_2_clka = io_clka; // @[util.scala 35:17]
  assign cluster_2_dina = io_dina; // @[util.scala 39:17]
  assign cluster_2_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_2_wea = io_wea & 18'h2 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_2_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_2_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_2_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_2_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_2_web = 1'h0; // @[util.scala 42:26]
  assign cluster_3_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_3_clka = io_clka; // @[util.scala 35:17]
  assign cluster_3_dina = io_dina; // @[util.scala 39:17]
  assign cluster_3_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_3_wea = io_wea & 18'h3 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_3_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_3_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_3_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_3_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_3_web = 1'h0; // @[util.scala 42:26]
  assign cluster_4_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_4_clka = io_clka; // @[util.scala 35:17]
  assign cluster_4_dina = io_dina; // @[util.scala 39:17]
  assign cluster_4_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_4_wea = io_wea & 18'h4 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_4_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_4_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_4_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_4_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_4_web = 1'h0; // @[util.scala 42:26]
  assign cluster_5_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_5_clka = io_clka; // @[util.scala 35:17]
  assign cluster_5_dina = io_dina; // @[util.scala 39:17]
  assign cluster_5_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_5_wea = io_wea & 18'h5 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_5_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_5_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_5_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_5_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_5_web = 1'h0; // @[util.scala 42:26]
  assign cluster_6_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_6_clka = io_clka; // @[util.scala 35:17]
  assign cluster_6_dina = io_dina; // @[util.scala 39:17]
  assign cluster_6_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_6_wea = io_wea & 18'h6 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_6_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_6_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_6_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_6_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_6_web = 1'h0; // @[util.scala 42:26]
  assign cluster_7_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_7_clka = io_clka; // @[util.scala 35:17]
  assign cluster_7_dina = io_dina; // @[util.scala 39:17]
  assign cluster_7_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_7_wea = io_wea & 18'h7 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_7_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_7_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_7_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_7_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_7_web = 1'h0; // @[util.scala 42:26]
  assign cluster_8_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_8_clka = io_clka; // @[util.scala 35:17]
  assign cluster_8_dina = io_dina; // @[util.scala 39:17]
  assign cluster_8_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_8_wea = io_wea & 18'h8 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_8_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_8_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_8_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_8_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_8_web = 1'h0; // @[util.scala 42:26]
  assign cluster_9_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_9_clka = io_clka; // @[util.scala 35:17]
  assign cluster_9_dina = io_dina; // @[util.scala 39:17]
  assign cluster_9_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_9_wea = io_wea & 18'h9 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_9_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_9_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_9_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_9_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_9_web = 1'h0; // @[util.scala 42:26]
  assign cluster_10_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_10_clka = io_clka; // @[util.scala 35:17]
  assign cluster_10_dina = io_dina; // @[util.scala 39:17]
  assign cluster_10_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_10_wea = io_wea & 18'ha == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_10_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_10_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_10_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_10_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_10_web = 1'h0; // @[util.scala 42:26]
  assign cluster_11_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_11_clka = io_clka; // @[util.scala 35:17]
  assign cluster_11_dina = io_dina; // @[util.scala 39:17]
  assign cluster_11_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_11_wea = io_wea & 18'hb == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_11_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_11_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_11_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_11_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_11_web = 1'h0; // @[util.scala 42:26]
  assign cluster_12_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_12_clka = io_clka; // @[util.scala 35:17]
  assign cluster_12_dina = io_dina; // @[util.scala 39:17]
  assign cluster_12_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_12_wea = io_wea & 18'hc == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_12_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_12_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_12_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_12_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_12_web = 1'h0; // @[util.scala 42:26]
  assign cluster_13_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_13_clka = io_clka; // @[util.scala 35:17]
  assign cluster_13_dina = io_dina; // @[util.scala 39:17]
  assign cluster_13_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_13_wea = io_wea & 18'hd == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_13_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_13_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_13_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_13_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_13_web = 1'h0; // @[util.scala 42:26]
  assign cluster_14_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_14_clka = io_clka; // @[util.scala 35:17]
  assign cluster_14_dina = io_dina; // @[util.scala 39:17]
  assign cluster_14_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_14_wea = io_wea & 18'he == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_14_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_14_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_14_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_14_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_14_web = 1'h0; // @[util.scala 42:26]
  assign cluster_15_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_15_clka = io_clka; // @[util.scala 35:17]
  assign cluster_15_dina = io_dina; // @[util.scala 39:17]
  assign cluster_15_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_15_wea = io_wea & 18'hf == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_15_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_15_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_15_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_15_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_15_web = 1'h0; // @[util.scala 42:26]
  assign cluster_16_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_16_clka = io_clka; // @[util.scala 35:17]
  assign cluster_16_dina = io_dina; // @[util.scala 39:17]
  assign cluster_16_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_16_wea = io_wea & 18'h10 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_16_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_16_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_16_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_16_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_16_web = 1'h0; // @[util.scala 42:26]
  assign cluster_17_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_17_clka = io_clka; // @[util.scala 35:17]
  assign cluster_17_dina = io_dina; // @[util.scala 39:17]
  assign cluster_17_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_17_wea = io_wea & 18'h11 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_17_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_17_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_17_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_17_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_17_web = 1'h0; // @[util.scala 42:26]
  assign cluster_18_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_18_clka = io_clka; // @[util.scala 35:17]
  assign cluster_18_dina = io_dina; // @[util.scala 39:17]
  assign cluster_18_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_18_wea = io_wea & 18'h12 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_18_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_18_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_18_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_18_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_18_web = 1'h0; // @[util.scala 42:26]
  assign cluster_19_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_19_clka = io_clka; // @[util.scala 35:17]
  assign cluster_19_dina = io_dina; // @[util.scala 39:17]
  assign cluster_19_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_19_wea = io_wea & 18'h13 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_19_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_19_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_19_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_19_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_19_web = 1'h0; // @[util.scala 42:26]
  assign cluster_20_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_20_clka = io_clka; // @[util.scala 35:17]
  assign cluster_20_dina = io_dina; // @[util.scala 39:17]
  assign cluster_20_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_20_wea = io_wea & 18'h14 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_20_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_20_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_20_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_20_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_20_web = 1'h0; // @[util.scala 42:26]
  assign cluster_21_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_21_clka = io_clka; // @[util.scala 35:17]
  assign cluster_21_dina = io_dina; // @[util.scala 39:17]
  assign cluster_21_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_21_wea = io_wea & 18'h15 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_21_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_21_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_21_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_21_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_21_web = 1'h0; // @[util.scala 42:26]
  assign cluster_22_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_22_clka = io_clka; // @[util.scala 35:17]
  assign cluster_22_dina = io_dina; // @[util.scala 39:17]
  assign cluster_22_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_22_wea = io_wea & 18'h16 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_22_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_22_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_22_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_22_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_22_web = 1'h0; // @[util.scala 42:26]
  assign cluster_23_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_23_clka = io_clka; // @[util.scala 35:17]
  assign cluster_23_dina = io_dina; // @[util.scala 39:17]
  assign cluster_23_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_23_wea = io_wea & 18'h17 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_23_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_23_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_23_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_23_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_23_web = 1'h0; // @[util.scala 42:26]
  assign cluster_24_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_24_clka = io_clka; // @[util.scala 35:17]
  assign cluster_24_dina = io_dina; // @[util.scala 39:17]
  assign cluster_24_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_24_wea = io_wea & 18'h18 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_24_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_24_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_24_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_24_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_24_web = 1'h0; // @[util.scala 42:26]
  assign cluster_25_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_25_clka = io_clka; // @[util.scala 35:17]
  assign cluster_25_dina = io_dina; // @[util.scala 39:17]
  assign cluster_25_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_25_wea = io_wea & 18'h19 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_25_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_25_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_25_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_25_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_25_web = 1'h0; // @[util.scala 42:26]
  assign cluster_26_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_26_clka = io_clka; // @[util.scala 35:17]
  assign cluster_26_dina = io_dina; // @[util.scala 39:17]
  assign cluster_26_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_26_wea = io_wea & 18'h1a == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_26_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_26_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_26_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_26_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_26_web = 1'h0; // @[util.scala 42:26]
  assign cluster_27_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_27_clka = io_clka; // @[util.scala 35:17]
  assign cluster_27_dina = io_dina; // @[util.scala 39:17]
  assign cluster_27_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_27_wea = io_wea & 18'h1b == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_27_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_27_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_27_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_27_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_27_web = 1'h0; // @[util.scala 42:26]
  assign cluster_28_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_28_clka = io_clka; // @[util.scala 35:17]
  assign cluster_28_dina = io_dina; // @[util.scala 39:17]
  assign cluster_28_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_28_wea = io_wea & 18'h1c == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_28_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_28_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_28_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_28_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_28_web = 1'h0; // @[util.scala 42:26]
  assign cluster_29_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_29_clka = io_clka; // @[util.scala 35:17]
  assign cluster_29_dina = io_dina; // @[util.scala 39:17]
  assign cluster_29_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_29_wea = io_wea & 18'h1d == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_29_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_29_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_29_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_29_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_29_web = 1'h0; // @[util.scala 42:26]
  assign cluster_30_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_30_clka = io_clka; // @[util.scala 35:17]
  assign cluster_30_dina = io_dina; // @[util.scala 39:17]
  assign cluster_30_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_30_wea = io_wea & 18'h1e == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_30_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_30_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_30_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_30_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_30_web = 1'h0; // @[util.scala 42:26]
  assign cluster_31_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_31_clka = io_clka; // @[util.scala 35:17]
  assign cluster_31_dina = io_dina; // @[util.scala 39:17]
  assign cluster_31_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_31_wea = io_wea & 18'h1f == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_31_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_31_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_31_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_31_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_31_web = 1'h0; // @[util.scala 42:26]
  assign cluster_32_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_32_clka = io_clka; // @[util.scala 35:17]
  assign cluster_32_dina = io_dina; // @[util.scala 39:17]
  assign cluster_32_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_32_wea = io_wea & 18'h20 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_32_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_32_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_32_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_32_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_32_web = 1'h0; // @[util.scala 42:26]
  assign cluster_33_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_33_clka = io_clka; // @[util.scala 35:17]
  assign cluster_33_dina = io_dina; // @[util.scala 39:17]
  assign cluster_33_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_33_wea = io_wea & 18'h21 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_33_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_33_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_33_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_33_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_33_web = 1'h0; // @[util.scala 42:26]
  assign cluster_34_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_34_clka = io_clka; // @[util.scala 35:17]
  assign cluster_34_dina = io_dina; // @[util.scala 39:17]
  assign cluster_34_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_34_wea = io_wea & 18'h22 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_34_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_34_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_34_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_34_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_34_web = 1'h0; // @[util.scala 42:26]
  assign cluster_35_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_35_clka = io_clka; // @[util.scala 35:17]
  assign cluster_35_dina = io_dina; // @[util.scala 39:17]
  assign cluster_35_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_35_wea = io_wea & 18'h23 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_35_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_35_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_35_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_35_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_35_web = 1'h0; // @[util.scala 42:26]
  assign cluster_36_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_36_clka = io_clka; // @[util.scala 35:17]
  assign cluster_36_dina = io_dina; // @[util.scala 39:17]
  assign cluster_36_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_36_wea = io_wea & 18'h24 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_36_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_36_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_36_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_36_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_36_web = 1'h0; // @[util.scala 42:26]
  assign cluster_37_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_37_clka = io_clka; // @[util.scala 35:17]
  assign cluster_37_dina = io_dina; // @[util.scala 39:17]
  assign cluster_37_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_37_wea = io_wea & 18'h25 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_37_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_37_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_37_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_37_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_37_web = 1'h0; // @[util.scala 42:26]
  assign cluster_38_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_38_clka = io_clka; // @[util.scala 35:17]
  assign cluster_38_dina = io_dina; // @[util.scala 39:17]
  assign cluster_38_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_38_wea = io_wea & 18'h26 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_38_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_38_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_38_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_38_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_38_web = 1'h0; // @[util.scala 42:26]
  assign cluster_39_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_39_clka = io_clka; // @[util.scala 35:17]
  assign cluster_39_dina = io_dina; // @[util.scala 39:17]
  assign cluster_39_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_39_wea = io_wea & 18'h27 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_39_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_39_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_39_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_39_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_39_web = 1'h0; // @[util.scala 42:26]
  assign cluster_40_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_40_clka = io_clka; // @[util.scala 35:17]
  assign cluster_40_dina = io_dina; // @[util.scala 39:17]
  assign cluster_40_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_40_wea = io_wea & 18'h28 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_40_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_40_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_40_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_40_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_40_web = 1'h0; // @[util.scala 42:26]
  assign cluster_41_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_41_clka = io_clka; // @[util.scala 35:17]
  assign cluster_41_dina = io_dina; // @[util.scala 39:17]
  assign cluster_41_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_41_wea = io_wea & 18'h29 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_41_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_41_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_41_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_41_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_41_web = 1'h0; // @[util.scala 42:26]
  assign cluster_42_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_42_clka = io_clka; // @[util.scala 35:17]
  assign cluster_42_dina = io_dina; // @[util.scala 39:17]
  assign cluster_42_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_42_wea = io_wea & 18'h2a == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_42_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_42_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_42_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_42_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_42_web = 1'h0; // @[util.scala 42:26]
  assign cluster_43_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_43_clka = io_clka; // @[util.scala 35:17]
  assign cluster_43_dina = io_dina; // @[util.scala 39:17]
  assign cluster_43_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_43_wea = io_wea & 18'h2b == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_43_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_43_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_43_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_43_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_43_web = 1'h0; // @[util.scala 42:26]
  assign cluster_44_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_44_clka = io_clka; // @[util.scala 35:17]
  assign cluster_44_dina = io_dina; // @[util.scala 39:17]
  assign cluster_44_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_44_wea = io_wea & 18'h2c == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_44_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_44_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_44_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_44_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_44_web = 1'h0; // @[util.scala 42:26]
  assign cluster_45_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_45_clka = io_clka; // @[util.scala 35:17]
  assign cluster_45_dina = io_dina; // @[util.scala 39:17]
  assign cluster_45_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_45_wea = io_wea & 18'h2d == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_45_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_45_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_45_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_45_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_45_web = 1'h0; // @[util.scala 42:26]
  assign cluster_46_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_46_clka = io_clka; // @[util.scala 35:17]
  assign cluster_46_dina = io_dina; // @[util.scala 39:17]
  assign cluster_46_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_46_wea = io_wea & 18'h2e == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_46_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_46_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_46_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_46_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_46_web = 1'h0; // @[util.scala 42:26]
  assign cluster_47_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_47_clka = io_clka; // @[util.scala 35:17]
  assign cluster_47_dina = io_dina; // @[util.scala 39:17]
  assign cluster_47_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_47_wea = io_wea & 18'h2f == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_47_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_47_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_47_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_47_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_47_web = 1'h0; // @[util.scala 42:26]
  assign cluster_48_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_48_clka = io_clka; // @[util.scala 35:17]
  assign cluster_48_dina = io_dina; // @[util.scala 39:17]
  assign cluster_48_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_48_wea = io_wea & 18'h30 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_48_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_48_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_48_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_48_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_48_web = 1'h0; // @[util.scala 42:26]
  assign cluster_49_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_49_clka = io_clka; // @[util.scala 35:17]
  assign cluster_49_dina = io_dina; // @[util.scala 39:17]
  assign cluster_49_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_49_wea = io_wea & 18'h31 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_49_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_49_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_49_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_49_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_49_web = 1'h0; // @[util.scala 42:26]
  assign cluster_50_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_50_clka = io_clka; // @[util.scala 35:17]
  assign cluster_50_dina = io_dina; // @[util.scala 39:17]
  assign cluster_50_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_50_wea = io_wea & 18'h32 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_50_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_50_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_50_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_50_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_50_web = 1'h0; // @[util.scala 42:26]
  assign cluster_51_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_51_clka = io_clka; // @[util.scala 35:17]
  assign cluster_51_dina = io_dina; // @[util.scala 39:17]
  assign cluster_51_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_51_wea = io_wea & 18'h33 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_51_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_51_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_51_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_51_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_51_web = 1'h0; // @[util.scala 42:26]
  assign cluster_52_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_52_clka = io_clka; // @[util.scala 35:17]
  assign cluster_52_dina = io_dina; // @[util.scala 39:17]
  assign cluster_52_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_52_wea = io_wea & 18'h34 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_52_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_52_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_52_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_52_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_52_web = 1'h0; // @[util.scala 42:26]
  assign cluster_53_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_53_clka = io_clka; // @[util.scala 35:17]
  assign cluster_53_dina = io_dina; // @[util.scala 39:17]
  assign cluster_53_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_53_wea = io_wea & 18'h35 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_53_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_53_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_53_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_53_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_53_web = 1'h0; // @[util.scala 42:26]
  assign cluster_54_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_54_clka = io_clka; // @[util.scala 35:17]
  assign cluster_54_dina = io_dina; // @[util.scala 39:17]
  assign cluster_54_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_54_wea = io_wea & 18'h36 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_54_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_54_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_54_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_54_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_54_web = 1'h0; // @[util.scala 42:26]
  assign cluster_55_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_55_clka = io_clka; // @[util.scala 35:17]
  assign cluster_55_dina = io_dina; // @[util.scala 39:17]
  assign cluster_55_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_55_wea = io_wea & 18'h37 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_55_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_55_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_55_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_55_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_55_web = 1'h0; // @[util.scala 42:26]
  assign cluster_56_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_56_clka = io_clka; // @[util.scala 35:17]
  assign cluster_56_dina = io_dina; // @[util.scala 39:17]
  assign cluster_56_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_56_wea = io_wea & 18'h38 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_56_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_56_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_56_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_56_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_56_web = 1'h0; // @[util.scala 42:26]
  assign cluster_57_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_57_clka = io_clka; // @[util.scala 35:17]
  assign cluster_57_dina = io_dina; // @[util.scala 39:17]
  assign cluster_57_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_57_wea = io_wea & 18'h39 == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_57_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_57_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_57_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_57_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_57_web = 1'h0; // @[util.scala 42:26]
  assign cluster_58_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_58_clka = io_clka; // @[util.scala 35:17]
  assign cluster_58_dina = io_dina; // @[util.scala 39:17]
  assign cluster_58_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_58_wea = io_wea & 18'h3a == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_58_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_58_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_58_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_58_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_58_web = 1'h0; // @[util.scala 42:26]
  assign cluster_59_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_59_clka = io_clka; // @[util.scala 35:17]
  assign cluster_59_dina = io_dina; // @[util.scala 39:17]
  assign cluster_59_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_59_wea = io_wea & 18'h3b == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_59_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_59_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_59_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_59_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_59_web = 1'h0; // @[util.scala 42:26]
  assign cluster_60_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_60_clka = io_clka; // @[util.scala 35:17]
  assign cluster_60_dina = io_dina; // @[util.scala 39:17]
  assign cluster_60_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_60_wea = io_wea & 18'h3c == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_60_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_60_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_60_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_60_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_60_web = 1'h0; // @[util.scala 42:26]
  assign cluster_61_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_61_clka = io_clka; // @[util.scala 35:17]
  assign cluster_61_dina = io_dina; // @[util.scala 39:17]
  assign cluster_61_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_61_wea = io_wea & 18'h3d == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_61_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_61_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_61_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_61_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_61_web = 1'h0; // @[util.scala 42:26]
  assign cluster_62_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_62_clka = io_clka; // @[util.scala 35:17]
  assign cluster_62_dina = io_dina; // @[util.scala 39:17]
  assign cluster_62_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_62_wea = io_wea & 18'h3e == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_62_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_62_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_62_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_62_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_62_web = 1'h0; // @[util.scala 42:26]
  assign cluster_63_addra = io_addra[11:0]; // @[util.scala 41:29]
  assign cluster_63_clka = io_clka; // @[util.scala 35:17]
  assign cluster_63_dina = io_dina; // @[util.scala 39:17]
  assign cluster_63_ena = 1'h1; // @[util.scala 37:16]
  assign cluster_63_wea = io_wea & 18'h3f == _cluster_0_io_wea_T; // @[util.scala 43:26]
  assign cluster_63_addrb = io_addrb[11:0]; // @[util.scala 40:29]
  assign cluster_63_clkb = io_clkb; // @[util.scala 34:17]
  assign cluster_63_dinb = 48'h0; // @[util.scala 38:17]
  assign cluster_63_enb = 1'h1; // @[util.scala 36:16]
  assign cluster_63_web = 1'h0; // @[util.scala 42:26]
endmodule
module pipeline_97(
  input         clock,
  input         reset,
  input         io_dout_ready,
  output        io_dout_valid,
  output [15:0] io_dout_bits_addr,
  output [11:0] io_dout_bits_block_index,
  output        io_din_ready,
  input         io_din_valid,
  input  [15:0] io_din_bits_addr,
  input  [11:0] io_din_bits_block_index
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] data_addr; // @[util.scala 143:21]
  reg [11:0] data_block_index; // @[util.scala 143:21]
  reg  valid; // @[util.scala 144:22]
  assign io_dout_valid = valid; // @[util.scala 151:17]
  assign io_dout_bits_addr = data_addr; // @[util.scala 152:16]
  assign io_dout_bits_block_index = data_block_index; // @[util.scala 152:16]
  assign io_din_ready = io_dout_ready; // @[util.scala 150:16]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 143:21]
      data_addr <= 16'h0; // @[util.scala 143:21]
    end else if (io_dout_ready) begin // @[util.scala 145:22]
      data_addr <= io_din_bits_addr; // @[util.scala 146:10]
    end
    if (reset) begin // @[util.scala 143:21]
      data_block_index <= 12'h0; // @[util.scala 143:21]
    end else if (io_dout_ready) begin // @[util.scala 145:22]
      data_block_index <= io_din_bits_block_index; // @[util.scala 146:10]
    end
    if (reset) begin // @[util.scala 144:22]
      valid <= 1'h0; // @[util.scala 144:22]
    end else if (io_dout_ready) begin // @[util.scala 145:22]
      valid <= io_din_valid; // @[util.scala 147:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_addr = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  data_block_index = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  valid = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WB_engine(
  input          clock,
  input          reset,
  input          io_ddr_aw_ready,
  output         io_ddr_aw_valid,
  output [63:0]  io_ddr_aw_bits_awaddr,
  output [6:0]   io_ddr_aw_bits_awid,
  input          io_ddr_w_ready,
  output         io_ddr_w_valid,
  output [511:0] io_ddr_w_bits_wdata,
  output [63:0]  io_ddr_w_bits_wstrb,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [31:0]  io_xbar_in_bits_tdata,
  input  [63:0]  io_level_base_addr,
  input  [31:0]  io_level,
  output         io_end,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [17:0] buffer_io_addra; // @[BFS.scala 24:22]
  wire  buffer_io_clka; // @[BFS.scala 24:22]
  wire [47:0] buffer_io_dina; // @[BFS.scala 24:22]
  wire  buffer_io_wea; // @[BFS.scala 24:22]
  wire [17:0] buffer_io_addrb; // @[BFS.scala 24:22]
  wire  buffer_io_clkb; // @[BFS.scala 24:22]
  wire [47:0] buffer_io_doutb; // @[BFS.scala 24:22]
  wire [11:0] region_counter__addra; // @[BFS.scala 25:30]
  wire  region_counter__clka; // @[BFS.scala 25:30]
  wire [8:0] region_counter__dina; // @[BFS.scala 25:30]
  wire  region_counter__ena; // @[BFS.scala 25:30]
  wire  region_counter__wea; // @[BFS.scala 25:30]
  wire [11:0] region_counter__addrb; // @[BFS.scala 25:30]
  wire  region_counter__clkb; // @[BFS.scala 25:30]
  wire [8:0] region_counter__doutb; // @[BFS.scala 25:30]
  wire  region_counter__enb; // @[BFS.scala 25:30]
  wire  region_counter_doutb_forward_clock; // @[BFS.scala 44:44]
  wire  region_counter_doutb_forward_reset; // @[BFS.scala 44:44]
  wire  region_counter_doutb_forward_io_dout_ready; // @[BFS.scala 44:44]
  wire  region_counter_doutb_forward_io_dout_valid; // @[BFS.scala 44:44]
  wire [8:0] region_counter_doutb_forward_io_dout_bits; // @[BFS.scala 44:44]
  wire  region_counter_doutb_forward_io_din_valid; // @[BFS.scala 44:44]
  wire [8:0] region_counter_doutb_forward_io_din_bits; // @[BFS.scala 44:44]
  wire  pipeline_1_clock; // @[BFS.scala 46:26]
  wire  pipeline_1_reset; // @[BFS.scala 46:26]
  wire  pipeline_1_io_dout_ready; // @[BFS.scala 46:26]
  wire  pipeline_1_io_dout_valid; // @[BFS.scala 46:26]
  wire [15:0] pipeline_1_io_dout_bits_addr; // @[BFS.scala 46:26]
  wire [11:0] pipeline_1_io_dout_bits_block_index; // @[BFS.scala 46:26]
  wire  pipeline_1_io_din_ready; // @[BFS.scala 46:26]
  wire  pipeline_1_io_din_valid; // @[BFS.scala 46:26]
  wire [15:0] pipeline_1_io_din_bits_addr; // @[BFS.scala 46:26]
  wire [11:0] pipeline_1_io_din_bits_block_index; // @[BFS.scala 46:26]
  wire  aw_buffer_full; // @[BFS.scala 79:25]
  wire [63:0] aw_buffer_din; // @[BFS.scala 79:25]
  wire  aw_buffer_wr_en; // @[BFS.scala 79:25]
  wire  aw_buffer_empty; // @[BFS.scala 79:25]
  wire [63:0] aw_buffer_dout; // @[BFS.scala 79:25]
  wire  aw_buffer_rd_en; // @[BFS.scala 79:25]
  wire [5:0] aw_buffer_data_count; // @[BFS.scala 79:25]
  wire  aw_buffer_clk; // @[BFS.scala 79:25]
  wire  aw_buffer_srst; // @[BFS.scala 79:25]
  wire  aw_buffer_valid; // @[BFS.scala 79:25]
  wire  w_buffer_full; // @[BFS.scala 80:24]
  wire [63:0] w_buffer_din; // @[BFS.scala 80:24]
  wire  w_buffer_wr_en; // @[BFS.scala 80:24]
  wire  w_buffer_empty; // @[BFS.scala 80:24]
  wire [63:0] w_buffer_dout; // @[BFS.scala 80:24]
  wire  w_buffer_rd_en; // @[BFS.scala 80:24]
  wire [5:0] w_buffer_data_count; // @[BFS.scala 80:24]
  wire  w_buffer_clk; // @[BFS.scala 80:24]
  wire  w_buffer_srst; // @[BFS.scala 80:24]
  wire  w_buffer_valid; // @[BFS.scala 80:24]
  wire [33:0] _GEN_16 = {io_xbar_in_bits_tdata, 2'h0}; // @[BFS.scala 34:23]
  wire [34:0] _dramaddr_T = {{1'd0}, _GEN_16}; // @[BFS.scala 34:23]
  wire [63:0] dramaddr = {{29'd0}, _dramaddr_T}; // @[BFS.scala 34:39 BFS.scala 34:39]
  wire [11:0] block_index = dramaddr[25:14]; // @[BFS.scala 35:29]
  wire  _pipeline_1_io_din_valid_T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 50:47]
  wire  _buffer_io_wea_T = pipeline_1_io_dout_valid & pipeline_1_io_dout_ready; // @[BFS.scala 56:45]
  wire [8:0] region_counter_doutb = region_counter_doutb_forward_io_dout_valid ?
    region_counter_doutb_forward_io_dout_bits : region_counter__doutb; // @[BFS.scala 68:30]
  wire [5:0] buffer_io_addra_lo = region_counter_doutb[5:0]; // @[BFS.scala 28:35 BFS.scala 28:35]
  wire [8:0] region_counter_dina_0 = region_counter_doutb + 9'h1; // @[BFS.scala 63:52]
  wire  _region_counter_doutb_forward_io_din_valid_T_1 = pipeline_1_io_dout_bits_block_index == block_index; // @[BFS.scala 66:28]
  wire  _region_counter_doutb_forward_io_din_valid_T_2 = _pipeline_1_io_din_valid_T &
    _region_counter_doutb_forward_io_din_valid_T_1; // @[BFS.scala 65:85]
  reg [1:0] wb_sm; // @[BFS.scala 77:22]
  reg [7:0] count; // @[BFS.scala 78:22]
  reg [11:0] wb_block_index; // @[BFS.scala 81:31]
  wire  _flush_start_T = wb_sm == 2'h0; // @[BFS.scala 82:28]
  wire  flush_start = wb_sm == 2'h0 & io_flush; // @[BFS.scala 82:42]
  reg [7:0] size_b; // @[BFS.scala 83:23]
  reg [63:0] level_base_addr_reg; // @[BFS.scala 84:36]
  wire  wb_start = pipeline_1_io_dout_valid & region_counter_doutb == 9'h3f; // @[BFS.scala 85:43]
  wire  _T = wb_sm == 2'h3; // @[BFS.scala 92:20]
  wire [8:0] _GEN_0 = wb_sm == 2'h3 ? region_counter_doutb : {{1'd0}, size_b}; // @[BFS.scala 92:38 BFS.scala 93:12 BFS.scala 83:23]
  wire [8:0] _GEN_1 = wb_start ? 9'h40 : _GEN_0; // @[BFS.scala 90:17 BFS.scala 91:12]
  wire  _T_1 = wb_sm == 2'h2; // @[BFS.scala 100:20]
  wire  _T_2 = wb_block_index != 12'hfff; // @[BFS.scala 100:55]
  wire [11:0] _wb_block_index_T_1 = wb_block_index + 12'h1; // @[BFS.scala 101:38]
  wire  _T_6 = wb_sm == 2'h1; // @[BFS.scala 115:20]
  wire  _T_7 = ~aw_buffer_full; // @[BFS.scala 115:57]
  wire  _T_9 = ~w_buffer_full; // @[BFS.scala 115:89]
  wire  _T_10 = wb_sm == 2'h1 & ~aw_buffer_full & ~w_buffer_full; // @[BFS.scala 115:69]
  wire [1:0] _GEN_6 = io_flush ? 2'h2 : 2'h0; // @[BFS.scala 117:21 BFS.scala 118:15 BFS.scala 120:15]
  wire [1:0] _GEN_7 = count == size_b ? _GEN_6 : 2'h1; // @[BFS.scala 116:27 BFS.scala 123:13]
  wire [1:0] _GEN_8 = _T_2 ? 2'h3 : 2'h0; // @[BFS.scala 126:46 BFS.scala 127:13 BFS.scala 129:13]
  wire [1:0] _GEN_9 = _T_1 ? _GEN_8 : wb_sm; // @[BFS.scala 125:38 BFS.scala 77:22]
  wire [1:0] _GEN_10 = wb_sm == 2'h1 & ~aw_buffer_full & ~w_buffer_full ? _GEN_7 : _GEN_9; // @[BFS.scala 115:102]
  wire [7:0] _count_T_1 = count + 8'h1; // @[BFS.scala 136:20]
  wire [17:0] _buffer_io_addrb_T = {block_index,6'h0}; // @[Cat.scala 30:58]
  wire [5:0] buffer_io_addrb_lo_2 = count[5:0]; // @[BFS.scala 28:35 BFS.scala 28:35]
  wire [17:0] _buffer_io_addrb_T_4 = {wb_block_index,buffer_io_addrb_lo_2}; // @[Cat.scala 30:58]
  wire [17:0] _buffer_io_addrb_T_5 = wb_start ? _buffer_io_addrb_T : 18'h0; // @[Mux.scala 27:72]
  wire [17:0] _buffer_io_addrb_T_6 = _T ? _buffer_io_addrb_T : 18'h0; // @[Mux.scala 27:72]
  wire [17:0] _buffer_io_addrb_T_7 = _T_6 ? _buffer_io_addrb_T_4 : 18'h0; // @[Mux.scala 27:72]
  wire [17:0] _buffer_io_addrb_T_8 = _buffer_io_addrb_T_5 | _buffer_io_addrb_T_6; // @[Mux.scala 27:72]
  wire [11:0] _region_counter_io_addrb_T_3 = flush_start ? 12'h0 : block_index; // @[Mux.scala 98:16]
  wire [13:0] aw_buffer_io_din_lo = buffer_io_doutb[45:32]; // @[BFS.scala 160:80]
  wire [25:0] _aw_buffer_io_din_T = {wb_block_index,aw_buffer_io_din_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_17 = {{38'd0}, _aw_buffer_io_din_T}; // @[BFS.scala 160:43]
  wire [57:0] alignment_addr = aw_buffer_dout[63:6]; // @[BFS.scala 161:41]
  wire [5:0] io_ddr_aw_bits_awid_lo = aw_buffer_data_count; // @[BFS.scala 164:72 BFS.scala 164:72]
  wire [5:0] alignment_offset = w_buffer_dout[37:32]; // @[BFS.scala 175:42]
  wire [9:0] _io_ddr_w_bits_wdata_T_1 = 4'h8 * alignment_offset; // @[BFS.scala 176:80]
  wire [511:0] _io_ddr_w_bits_wdata_WIRE = {{480'd0}, w_buffer_dout[31:0]}; // @[BFS.scala 176:58 BFS.scala 176:58]
  wire [1534:0] _GEN_18 = {{1023'd0}, _io_ddr_w_bits_wdata_WIRE}; // @[BFS.scala 176:72]
  wire [1534:0] _io_ddr_w_bits_wdata_T_2 = _GEN_18 << _io_ddr_w_bits_wdata_T_1; // @[BFS.scala 176:72]
  wire [126:0] _io_ddr_w_bits_wstrb_T = 127'hf << alignment_offset; // @[BFS.scala 179:38]
  URAM_cluster buffer ( // @[BFS.scala 24:22]
    .io_addra(buffer_io_addra),
    .io_clka(buffer_io_clka),
    .io_dina(buffer_io_dina),
    .io_wea(buffer_io_wea),
    .io_addrb(buffer_io_addrb),
    .io_clkb(buffer_io_clkb),
    .io_doutb(buffer_io_doutb)
  );
  region_counter region_counter_ ( // @[BFS.scala 25:30]
    .addra(region_counter__addra),
    .clka(region_counter__clka),
    .dina(region_counter__dina),
    .ena(region_counter__ena),
    .wea(region_counter__wea),
    .addrb(region_counter__addrb),
    .clkb(region_counter__clkb),
    .doutb(region_counter__doutb),
    .enb(region_counter__enb)
  );
  pipeline_34 region_counter_doutb_forward ( // @[BFS.scala 44:44]
    .clock(region_counter_doutb_forward_clock),
    .reset(region_counter_doutb_forward_reset),
    .io_dout_ready(region_counter_doutb_forward_io_dout_ready),
    .io_dout_valid(region_counter_doutb_forward_io_dout_valid),
    .io_dout_bits(region_counter_doutb_forward_io_dout_bits),
    .io_din_valid(region_counter_doutb_forward_io_din_valid),
    .io_din_bits(region_counter_doutb_forward_io_din_bits)
  );
  pipeline_97 pipeline_1 ( // @[BFS.scala 46:26]
    .clock(pipeline_1_clock),
    .reset(pipeline_1_reset),
    .io_dout_ready(pipeline_1_io_dout_ready),
    .io_dout_valid(pipeline_1_io_dout_valid),
    .io_dout_bits_addr(pipeline_1_io_dout_bits_addr),
    .io_dout_bits_block_index(pipeline_1_io_dout_bits_block_index),
    .io_din_ready(pipeline_1_io_din_ready),
    .io_din_valid(pipeline_1_io_din_valid),
    .io_din_bits_addr(pipeline_1_io_din_bits_addr),
    .io_din_bits_block_index(pipeline_1_io_din_bits_block_index)
  );
  addr_fifo aw_buffer ( // @[BFS.scala 79:25]
    .full(aw_buffer_full),
    .din(aw_buffer_din),
    .wr_en(aw_buffer_wr_en),
    .empty(aw_buffer_empty),
    .dout(aw_buffer_dout),
    .rd_en(aw_buffer_rd_en),
    .data_count(aw_buffer_data_count),
    .clk(aw_buffer_clk),
    .srst(aw_buffer_srst),
    .valid(aw_buffer_valid)
  );
  level_fifo w_buffer ( // @[BFS.scala 80:24]
    .full(w_buffer_full),
    .din(w_buffer_din),
    .wr_en(w_buffer_wr_en),
    .empty(w_buffer_empty),
    .dout(w_buffer_dout),
    .rd_en(w_buffer_rd_en),
    .data_count(w_buffer_data_count),
    .clk(w_buffer_clk),
    .srst(w_buffer_srst),
    .valid(w_buffer_valid)
  );
  assign io_ddr_aw_valid = aw_buffer_valid; // @[BFS.scala 168:19]
  assign io_ddr_aw_bits_awaddr = {alignment_addr,6'h0}; // @[Cat.scala 30:58]
  assign io_ddr_aw_bits_awid = {1'h1,io_ddr_aw_bits_awid_lo}; // @[Cat.scala 30:58]
  assign io_ddr_w_valid = w_buffer_valid; // @[BFS.scala 178:18]
  assign io_ddr_w_bits_wdata = _io_ddr_w_bits_wdata_T_2[511:0]; // @[BFS.scala 176:23]
  assign io_ddr_w_bits_wstrb = _io_ddr_w_bits_wstrb_T[63:0]; // @[BFS.scala 179:23]
  assign io_xbar_in_ready = pipeline_1_io_din_ready; // @[BFS.scala 53:20]
  assign io_end = _T_1 & wb_block_index == 12'hfff; // @[BFS.scala 184:36]
  assign buffer_io_addra = {pipeline_1_io_dout_bits_block_index,buffer_io_addra_lo}; // @[Cat.scala 30:58]
  assign buffer_io_clka = clock; // @[BFS.scala 59:33]
  assign buffer_io_dina = {pipeline_1_io_dout_bits_addr,io_level}; // @[Cat.scala 30:58]
  assign buffer_io_wea = pipeline_1_io_dout_valid & pipeline_1_io_dout_ready; // @[BFS.scala 56:45]
  assign buffer_io_addrb = _buffer_io_addrb_T_8 | _buffer_io_addrb_T_7; // @[Mux.scala 27:72]
  assign buffer_io_clkb = clock; // @[BFS.scala 147:33]
  assign region_counter__addra = _T_6 ? wb_block_index : pipeline_1_io_dout_bits_block_index; // @[BFS.scala 149:33]
  assign region_counter__clka = clock; // @[BFS.scala 38:41]
  assign region_counter__dina = _T_6 ? 9'h0 : region_counter_dina_0; // @[BFS.scala 151:32]
  assign region_counter__ena = 1'h1; // @[BFS.scala 39:25]
  assign region_counter__wea = _T_6 | _buffer_io_wea_T; // @[BFS.scala 150:31]
  assign region_counter__addrb = _T_1 ? _wb_block_index_T_1 : _region_counter_io_addrb_T_3; // @[Mux.scala 98:16]
  assign region_counter__clkb = clock; // @[BFS.scala 37:41]
  assign region_counter__enb = 1'h1; // @[BFS.scala 40:25]
  assign region_counter_doutb_forward_clock = clock;
  assign region_counter_doutb_forward_reset = reset;
  assign region_counter_doutb_forward_io_dout_ready = wb_sm == 2'h0; // @[BFS.scala 87:55]
  assign region_counter_doutb_forward_io_din_valid = _region_counter_doutb_forward_io_din_valid_T_2 & _buffer_io_wea_T; // @[BFS.scala 66:55]
  assign region_counter_doutb_forward_io_din_bits = region_counter_doutb + 9'h1; // @[BFS.scala 63:52]
  assign pipeline_1_clock = clock;
  assign pipeline_1_reset = reset;
  assign pipeline_1_io_dout_ready = wb_sm == 2'h0; // @[BFS.scala 86:37]
  assign pipeline_1_io_din_valid = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 50:47]
  assign pipeline_1_io_din_bits_addr = {{2'd0}, dramaddr[13:0]}; // @[BFS.scala 51:58 BFS.scala 51:58]
  assign pipeline_1_io_din_bits_block_index = dramaddr[25:14]; // @[BFS.scala 35:29]
  assign aw_buffer_din = level_base_addr_reg + _GEN_17; // @[BFS.scala 160:43]
  assign aw_buffer_wr_en = _T_6 & _T_9; // @[BFS.scala 159:47]
  assign aw_buffer_rd_en = io_ddr_aw_ready; // @[BFS.scala 169:22]
  assign aw_buffer_clk = clock; // @[BFS.scala 157:35]
  assign aw_buffer_srst = reset; // @[BFS.scala 158:36]
  assign w_buffer_din = {{26'd0}, buffer_io_doutb[37:0]}; // @[BFS.scala 174:37]
  assign w_buffer_wr_en = _T_6 & _T_7; // @[BFS.scala 173:46]
  assign w_buffer_rd_en = io_ddr_w_ready; // @[BFS.scala 180:21]
  assign w_buffer_clk = clock; // @[BFS.scala 171:34]
  assign w_buffer_srst = reset; // @[BFS.scala 172:35]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 77:22]
      wb_sm <= 2'h0; // @[BFS.scala 77:22]
    end else if (flush_start) begin // @[BFS.scala 105:20]
      wb_sm <= 2'h3; // @[BFS.scala 106:11]
    end else if (_T) begin // @[BFS.scala 107:38]
      if (region_counter_doutb == 9'h0) begin // @[BFS.scala 108:39]
        wb_sm <= 2'h2; // @[BFS.scala 109:13]
      end else begin
        wb_sm <= 2'h1; // @[BFS.scala 111:13]
      end
    end else if (wb_start) begin // @[BFS.scala 113:23]
      wb_sm <= 2'h1; // @[BFS.scala 114:11]
    end else begin
      wb_sm <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 78:22]
      count <= 8'h0; // @[BFS.scala 78:22]
    end else if (_flush_start_T | _T_1) begin // @[BFS.scala 133:53]
      count <= 8'h1; // @[BFS.scala 134:11]
    end else if (_T_10) begin // @[BFS.scala 135:101]
      count <= _count_T_1; // @[BFS.scala 136:11]
    end
    if (reset) begin // @[BFS.scala 81:31]
      wb_block_index <= 12'h0; // @[BFS.scala 81:31]
    end else if (wb_start) begin // @[BFS.scala 96:17]
      wb_block_index <= pipeline_1_io_dout_bits_block_index; // @[BFS.scala 97:20]
    end else if (flush_start) begin // @[BFS.scala 98:26]
      wb_block_index <= 12'h0; // @[BFS.scala 99:20]
    end else if (wb_sm == 2'h2 & wb_block_index != 12'hfff) begin // @[BFS.scala 100:76]
      wb_block_index <= _wb_block_index_T_1; // @[BFS.scala 101:20]
    end
    if (reset) begin // @[BFS.scala 83:23]
      size_b <= 8'h0; // @[BFS.scala 83:23]
    end else begin
      size_b <= _GEN_1[7:0];
    end
    if (reset) begin // @[BFS.scala 84:36]
      level_base_addr_reg <= 64'h0; // @[BFS.scala 84:36]
    end else begin
      level_base_addr_reg <= io_level_base_addr; // @[BFS.scala 88:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_sm = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  wb_block_index = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  size_b = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  level_base_addr_reg = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Apply(
  input          clock,
  input          reset,
  input          io_ddr_aw_ready,
  output         io_ddr_aw_valid,
  output [63:0]  io_ddr_aw_bits_awaddr,
  output [6:0]   io_ddr_aw_bits_awid,
  input          io_ddr_w_ready,
  output         io_ddr_w_valid,
  output [511:0] io_ddr_w_bits_wdata,
  output [63:0]  io_ddr_w_bits_wstrb,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input  [31:0]  io_level,
  input  [63:0]  io_level_base_addr,
  output         io_end,
  input          io_flush
);
  wire  vertex_update_buffer_full; // @[BFS.scala 204:36]
  wire [63:0] vertex_update_buffer_din; // @[BFS.scala 204:36]
  wire  vertex_update_buffer_wr_en; // @[BFS.scala 204:36]
  wire  vertex_update_buffer_empty; // @[BFS.scala 204:36]
  wire [63:0] vertex_update_buffer_dout; // @[BFS.scala 204:36]
  wire  vertex_update_buffer_rd_en; // @[BFS.scala 204:36]
  wire [5:0] vertex_update_buffer_data_count; // @[BFS.scala 204:36]
  wire  vertex_update_buffer_clk; // @[BFS.scala 204:36]
  wire  vertex_update_buffer_srst; // @[BFS.scala 204:36]
  wire  vertex_update_buffer_valid; // @[BFS.scala 204:36]
  wire  update_engine_clock; // @[BFS.scala 213:29]
  wire  update_engine_reset; // @[BFS.scala 213:29]
  wire  update_engine_io_ddr_aw_ready; // @[BFS.scala 213:29]
  wire  update_engine_io_ddr_aw_valid; // @[BFS.scala 213:29]
  wire [63:0] update_engine_io_ddr_aw_bits_awaddr; // @[BFS.scala 213:29]
  wire [6:0] update_engine_io_ddr_aw_bits_awid; // @[BFS.scala 213:29]
  wire  update_engine_io_ddr_w_ready; // @[BFS.scala 213:29]
  wire  update_engine_io_ddr_w_valid; // @[BFS.scala 213:29]
  wire [511:0] update_engine_io_ddr_w_bits_wdata; // @[BFS.scala 213:29]
  wire [63:0] update_engine_io_ddr_w_bits_wstrb; // @[BFS.scala 213:29]
  wire  update_engine_io_xbar_in_ready; // @[BFS.scala 213:29]
  wire  update_engine_io_xbar_in_valid; // @[BFS.scala 213:29]
  wire [31:0] update_engine_io_xbar_in_bits_tdata; // @[BFS.scala 213:29]
  wire [63:0] update_engine_io_level_base_addr; // @[BFS.scala 213:29]
  wire [31:0] update_engine_io_level; // @[BFS.scala 213:29]
  wire  update_engine_io_end; // @[BFS.scala 213:29]
  wire  update_engine_io_flush; // @[BFS.scala 213:29]
  wire  FIN = io_gather_in_bits_tdata[31] & io_gather_in_valid; // @[BFS.scala 205:41]
  wire  _update_engine_io_flush_T = vertex_update_buffer_data_count == 6'h0; // @[util.scala 116:19]
  update_fifo vertex_update_buffer ( // @[BFS.scala 204:36]
    .full(vertex_update_buffer_full),
    .din(vertex_update_buffer_din),
    .wr_en(vertex_update_buffer_wr_en),
    .empty(vertex_update_buffer_empty),
    .dout(vertex_update_buffer_dout),
    .rd_en(vertex_update_buffer_rd_en),
    .data_count(vertex_update_buffer_data_count),
    .clk(vertex_update_buffer_clk),
    .srst(vertex_update_buffer_srst),
    .valid(vertex_update_buffer_valid)
  );
  WB_engine update_engine ( // @[BFS.scala 213:29]
    .clock(update_engine_clock),
    .reset(update_engine_reset),
    .io_ddr_aw_ready(update_engine_io_ddr_aw_ready),
    .io_ddr_aw_valid(update_engine_io_ddr_aw_valid),
    .io_ddr_aw_bits_awaddr(update_engine_io_ddr_aw_bits_awaddr),
    .io_ddr_aw_bits_awid(update_engine_io_ddr_aw_bits_awid),
    .io_ddr_w_ready(update_engine_io_ddr_w_ready),
    .io_ddr_w_valid(update_engine_io_ddr_w_valid),
    .io_ddr_w_bits_wdata(update_engine_io_ddr_w_bits_wdata),
    .io_ddr_w_bits_wstrb(update_engine_io_ddr_w_bits_wstrb),
    .io_xbar_in_ready(update_engine_io_xbar_in_ready),
    .io_xbar_in_valid(update_engine_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(update_engine_io_xbar_in_bits_tdata),
    .io_level_base_addr(update_engine_io_level_base_addr),
    .io_level(update_engine_io_level),
    .io_end(update_engine_io_end),
    .io_flush(update_engine_io_flush)
  );
  assign io_ddr_aw_valid = update_engine_io_ddr_aw_valid; // @[BFS.scala 223:13]
  assign io_ddr_aw_bits_awaddr = update_engine_io_ddr_aw_bits_awaddr; // @[BFS.scala 223:13]
  assign io_ddr_aw_bits_awid = update_engine_io_ddr_aw_bits_awid; // @[BFS.scala 223:13]
  assign io_ddr_w_valid = update_engine_io_ddr_w_valid; // @[BFS.scala 224:12]
  assign io_ddr_w_bits_wdata = update_engine_io_ddr_w_bits_wdata; // @[BFS.scala 224:12]
  assign io_ddr_w_bits_wstrb = update_engine_io_ddr_w_bits_wstrb; // @[BFS.scala 224:12]
  assign io_gather_in_ready = ~vertex_update_buffer_full; // @[BFS.scala 211:54]
  assign io_end = update_engine_io_end; // @[BFS.scala 226:10]
  assign vertex_update_buffer_din = {io_gather_in_bits_tdata,io_level}; // @[Cat.scala 30:58]
  assign vertex_update_buffer_wr_en = io_gather_in_valid & ~FIN; // @[BFS.scala 208:55]
  assign vertex_update_buffer_rd_en = update_engine_io_xbar_in_ready; // @[BFS.scala 221:33]
  assign vertex_update_buffer_clk = clock; // @[BFS.scala 206:46]
  assign vertex_update_buffer_srst = reset; // @[BFS.scala 207:47]
  assign update_engine_clock = clock;
  assign update_engine_reset = reset;
  assign update_engine_io_ddr_aw_ready = io_ddr_aw_ready; // @[BFS.scala 223:13]
  assign update_engine_io_ddr_w_ready = io_ddr_w_ready; // @[BFS.scala 224:12]
  assign update_engine_io_xbar_in_valid = vertex_update_buffer_valid; // @[BFS.scala 215:34]
  assign update_engine_io_xbar_in_bits_tdata = vertex_update_buffer_dout[63:32]; // @[BFS.scala 214:70]
  assign update_engine_io_level_base_addr = io_level_base_addr; // @[BFS.scala 216:36]
  assign update_engine_io_level = vertex_update_buffer_dout[31:0]; // @[BFS.scala 220:57]
  assign update_engine_io_flush = io_flush & _update_engine_io_flush_T; // @[BFS.scala 227:38]
endmodule
module readEdge_engine(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_rdata,
  input  [5:0]   io_in_bits_rid,
  input          io_in_bits_rlast,
  input          io_out_ready,
  output         io_out_valid,
  output [63:0]  io_out_bits_araddr,
  output [5:0]   io_out_bits_arid,
  output [7:0]   io_out_bits_arlen,
  output [2:0]   io_out_bits_arsize,
  input  [63:0]  io_edge_base_addr,
  input  [4:0]   io_free_ptr,
  output [31:0]  io_read_edge_num
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  edge_read_buffer_full; // @[BFS.scala 369:32]
  wire [63:0] edge_read_buffer_din; // @[BFS.scala 369:32]
  wire  edge_read_buffer_wr_en; // @[BFS.scala 369:32]
  wire  edge_read_buffer_empty; // @[BFS.scala 369:32]
  wire [63:0] edge_read_buffer_dout; // @[BFS.scala 369:32]
  wire  edge_read_buffer_rd_en; // @[BFS.scala 369:32]
  wire [5:0] edge_read_buffer_data_count; // @[BFS.scala 369:32]
  wire  edge_read_buffer_clk; // @[BFS.scala 369:32]
  wire  edge_read_buffer_srst; // @[BFS.scala 369:32]
  wire  edge_read_buffer_valid; // @[BFS.scala 369:32]
  reg  transaction_start; // @[BFS.scala 370:34]
  wire  _T = io_in_valid & io_in_ready; // @[BFS.scala 371:20]
  wire  _GEN_0 = _T & io_in_bits_rlast ? 1'h0 : transaction_start; // @[BFS.scala 373:70 BFS.scala 374:23 BFS.scala 370:34]
  wire  _GEN_1 = io_in_valid & io_in_ready & ~io_in_bits_rlast | _GEN_0; // @[BFS.scala 371:66 BFS.scala 372:23]
  wire  _edge_read_buffer_io_wr_en_T_5 = io_in_bits_rdata[63:32] > 32'he; // @[BFS.scala 380:39]
  wire  _edge_read_buffer_io_wr_en_T_6 = ~io_in_bits_rid[5] & io_in_valid & _edge_read_buffer_io_wr_en_T_5; // @[BFS.scala 379:72]
  wire [31:0] remainning_edges = edge_read_buffer_dout[63:32] - 32'he; // @[BFS.scala 383:68]
  reg  cache_status; // @[BFS.scala 389:29]
  reg [31:0] counter; // @[BFS.scala 390:24]
  reg [63:0] araddr; // @[BFS.scala 392:23]
  wire [31:0] next_counter = counter - 32'h40; // @[BFS.scala 394:27]
  wire  _T_10 = ~cache_status; // @[BFS.scala 395:116]
  wire [31:0] _counter_T_1 = remainning_edges - 32'h40; // @[BFS.scala 397:33]
  wire [33:0] _araddr_T_1 = {edge_read_buffer_dout[31:0], 2'h0}; // @[BFS.scala 398:83]
  wire [63:0] _GEN_11 = {{30'd0}, _araddr_T_1}; // @[BFS.scala 398:33]
  wire [63:0] _araddr_T_3 = io_edge_base_addr + _GEN_11; // @[BFS.scala 398:33]
  wire [63:0] _araddr_T_6 = _araddr_T_3 + 64'h100; // @[BFS.scala 398:98]
  wire  _T_15 = counter <= 32'h40; // @[BFS.scala 400:18]
  wire [63:0] _araddr_T_9 = araddr + 64'h100; // @[BFS.scala 406:24]
  wire  _GEN_2 = counter <= 32'h40 ? 1'h0 : cache_status; // @[BFS.scala 400:53 BFS.scala 401:20 BFS.scala 389:29]
  wire  _GEN_5 = io_out_ready & io_out_valid & cache_status ? _GEN_2 : cache_status; // @[BFS.scala 399:82 BFS.scala 389:29]
  wire  _GEN_8 = remainning_edges > 32'h40 & io_out_ready & io_out_valid & ~cache_status | _GEN_5; // @[BFS.scala 395:135 BFS.scala 396:18]
  wire  _num_vertex_T_2 = _T_10 & remainning_edges <= 32'h40; // @[BFS.scala 411:38]
  wire  _num_vertex_T_5 = cache_status & _T_15; // @[BFS.scala 412:42]
  wire [31:0] _num_vertex_T_6 = _num_vertex_T_5 ? counter : 32'h40; // @[Mux.scala 98:16]
  wire [31:0] num_vertex = _num_vertex_T_2 ? remainning_edges : _num_vertex_T_6; // @[Mux.scala 98:16]
  wire [31:0] _arlen_T_1 = {num_vertex[31:2], 2'h0}; // @[BFS.scala 414:63]
  wire [29:0] _arlen_T_6 = num_vertex[31:2] - 30'h1; // @[BFS.scala 416:57]
  wire [29:0] arlen = _arlen_T_1 < num_vertex ? num_vertex[31:2] : _arlen_T_6; // @[BFS.scala 414:18]
  wire  _io_out_bits_arsize_T = num_vertex <= 32'h1; // @[BFS.scala 425:23]
  wire  _io_out_bits_arsize_T_1 = num_vertex <= 32'h2; // @[BFS.scala 425:23]
  wire [2:0] _io_out_bits_arsize_T_2 = _io_out_bits_arsize_T_1 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  meta_fifo edge_read_buffer ( // @[BFS.scala 369:32]
    .full(edge_read_buffer_full),
    .din(edge_read_buffer_din),
    .wr_en(edge_read_buffer_wr_en),
    .empty(edge_read_buffer_empty),
    .dout(edge_read_buffer_dout),
    .rd_en(edge_read_buffer_rd_en),
    .data_count(edge_read_buffer_data_count),
    .clk(edge_read_buffer_clk),
    .srst(edge_read_buffer_srst),
    .valid(edge_read_buffer_valid)
  );
  assign io_in_ready = ~edge_read_buffer_full; // @[BFS.scala 381:43]
  assign io_out_valid = _T_10 ? edge_read_buffer_valid : 1'h1; // @[BFS.scala 420:22]
  assign io_out_bits_araddr = _T_10 ? _araddr_T_3 : araddr; // @[BFS.scala 417:28]
  assign io_out_bits_arid = {1'h1,io_free_ptr}; // @[Cat.scala 30:58]
  assign io_out_bits_arlen = arlen[7:0]; // @[BFS.scala 421:21]
  assign io_out_bits_arsize = _io_out_bits_arsize_T ? 3'h2 : _io_out_bits_arsize_T_2; // @[Mux.scala 98:16]
  assign io_read_edge_num = _num_vertex_T_2 ? remainning_edges : _num_vertex_T_6; // @[Mux.scala 98:16]
  assign edge_read_buffer_din = io_in_bits_rdata[63:0]; // @[BFS.scala 378:46]
  assign edge_read_buffer_wr_en = _edge_read_buffer_io_wr_en_T_6 & ~transaction_start; // @[BFS.scala 380:61]
  assign edge_read_buffer_rd_en = io_out_ready & _T_10; // @[BFS.scala 434:45]
  assign edge_read_buffer_clk = clock; // @[BFS.scala 376:42]
  assign edge_read_buffer_srst = reset; // @[BFS.scala 377:43]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 370:34]
      transaction_start <= 1'h0; // @[BFS.scala 370:34]
    end else begin
      transaction_start <= _GEN_1;
    end
    if (reset) begin // @[BFS.scala 389:29]
      cache_status <= 1'h0; // @[BFS.scala 389:29]
    end else begin
      cache_status <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 390:24]
      counter <= 32'h0; // @[BFS.scala 390:24]
    end else if (remainning_edges > 32'h40 & io_out_ready & io_out_valid & ~cache_status) begin // @[BFS.scala 395:135]
      counter <= _counter_T_1; // @[BFS.scala 397:13]
    end else if (io_out_ready & io_out_valid & cache_status) begin // @[BFS.scala 399:82]
      if (counter <= 32'h40) begin // @[BFS.scala 400:53]
        counter <= 32'h0; // @[BFS.scala 402:15]
      end else begin
        counter <= next_counter; // @[BFS.scala 405:15]
      end
    end
    if (reset) begin // @[BFS.scala 392:23]
      araddr <= 64'h0; // @[BFS.scala 392:23]
    end else if (remainning_edges > 32'h40 & io_out_ready & io_out_valid & ~cache_status) begin // @[BFS.scala 395:135]
      araddr <= _araddr_T_6; // @[BFS.scala 398:12]
    end else if (io_out_ready & io_out_valid & cache_status) begin // @[BFS.scala 399:82]
      if (counter <= 32'h40) begin // @[BFS.scala 400:53]
        araddr <= 64'h0; // @[BFS.scala 403:14]
      end else begin
        araddr <= _araddr_T_9; // @[BFS.scala 406:14]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  transaction_start = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cache_status = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  araddr = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AMBA_Arbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_araddr,
  input  [5:0]  io_in_0_bits_arid,
  input  [7:0]  io_in_0_bits_arlen,
  input  [2:0]  io_in_0_bits_arsize,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_araddr,
  input  [5:0]  io_in_1_bits_arid,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_araddr,
  output [5:0]  io_out_bits_arid,
  output [7:0]  io_out_bits_arlen,
  output [2:0]  io_out_bits_arsize
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  status; // @[util.scala 206:23]
  wire  grant_1 = ~io_in_0_valid; // @[util.scala 195:78]
  reg  grant_reg_0; // @[util.scala 208:26]
  reg  grant_reg_1; // @[util.scala 208:26]
  wire  _T = ~status; // @[util.scala 213:17]
  wire [2:0] _GEN_3 = io_in_0_valid ? io_in_0_bits_arsize : 3'h4; // @[util.scala 214:28 util.scala 216:21 util.scala 211:15]
  wire [7:0] _GEN_4 = io_in_0_valid ? io_in_0_bits_arlen : 8'h3; // @[util.scala 214:28 util.scala 216:21 util.scala 211:15]
  wire [5:0] _GEN_5 = io_in_0_valid ? io_in_0_bits_arid : io_in_1_bits_arid; // @[util.scala 214:28 util.scala 216:21 util.scala 211:15]
  wire [63:0] _GEN_6 = io_in_0_valid ? io_in_0_bits_araddr : io_in_1_bits_araddr; // @[util.scala 214:28 util.scala 216:21 util.scala 211:15]
  wire [2:0] _GEN_10 = grant_reg_0 ? io_in_0_bits_arsize : 3'h4; // @[util.scala 219:26 util.scala 221:21 util.scala 211:15]
  wire [7:0] _GEN_11 = grant_reg_0 ? io_in_0_bits_arlen : 8'h3; // @[util.scala 219:26 util.scala 221:21 util.scala 211:15]
  wire [5:0] _GEN_12 = grant_reg_0 ? io_in_0_bits_arid : io_in_1_bits_arid; // @[util.scala 219:26 util.scala 221:21 util.scala 211:15]
  wire [63:0] _GEN_13 = grant_reg_0 ? io_in_0_bits_araddr : io_in_1_bits_araddr; // @[util.scala 219:26 util.scala 221:21 util.scala 211:15]
  wire [2:0] _GEN_17 = status ? _GEN_10 : 3'h4; // @[util.scala 218:35 util.scala 211:15]
  wire [7:0] _GEN_18 = status ? _GEN_11 : 8'h3; // @[util.scala 218:35 util.scala 211:15]
  wire [5:0] _GEN_19 = status ? _GEN_12 : io_in_1_bits_arid; // @[util.scala 218:35 util.scala 211:15]
  wire [63:0] _GEN_20 = status ? _GEN_13 : io_in_1_bits_araddr; // @[util.scala 218:35 util.scala 211:15]
  wire  _T_6 = grant_1 & io_in_1_valid; // @[util.scala 228:24]
  wire  _GEN_28 = io_out_valid & io_out_ready & status ? 1'h0 : status; // @[util.scala 231:66 util.scala 232:12 util.scala 206:23]
  wire  _GEN_31 = (io_in_0_valid | io_in_1_valid) & _T | _GEN_28; // @[util.scala 226:62 util.scala 230:12]
  assign io_in_0_ready = _T ? io_out_ready : grant_reg_0 & io_out_ready; // @[util.scala 235:20]
  assign io_in_1_ready = _T ? grant_1 & io_out_ready : grant_reg_1 & io_out_ready; // @[util.scala 235:20]
  assign io_out_valid = _T ? ~grant_1 | io_in_1_valid : ~grant_reg_1 | io_in_1_valid; // @[util.scala 237:22]
  assign io_out_bits_araddr = ~status ? _GEN_6 : _GEN_20; // @[util.scala 213:30]
  assign io_out_bits_arid = ~status ? _GEN_5 : _GEN_19; // @[util.scala 213:30]
  assign io_out_bits_arlen = ~status ? _GEN_4 : _GEN_18; // @[util.scala 213:30]
  assign io_out_bits_arsize = ~status ? _GEN_3 : _GEN_17; // @[util.scala 213:30]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 206:23]
      status <= 1'h0; // @[util.scala 206:23]
    end else begin
      status <= _GEN_31;
    end
    if (reset) begin // @[util.scala 208:26]
      grant_reg_0 <= 1'h0; // @[util.scala 208:26]
    end else if ((io_in_0_valid | io_in_1_valid) & _T) begin // @[util.scala 226:62]
      grant_reg_0 <= io_in_0_valid; // @[util.scala 227:15]
    end
    if (reset) begin // @[util.scala 208:26]
      grant_reg_1 <= 1'h0; // @[util.scala 208:26]
    end else if ((io_in_0_valid | io_in_1_valid) & _T) begin // @[util.scala 226:62]
      grant_reg_1 <= _T_6; // @[util.scala 227:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  status = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  grant_reg_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  grant_reg_1 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module regFile(
  input         clock,
  input         reset,
  input  [31:0] io_dataIn,
  output [31:0] io_dataOut,
  input         io_writeFlag,
  input  [4:0]  io_rptr,
  input  [4:0]  io_wptr,
  output [4:0]  io_wcount
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[util.scala 83:21]
  reg [31:0] regs_1; // @[util.scala 83:21]
  reg [31:0] regs_2; // @[util.scala 83:21]
  reg [31:0] regs_3; // @[util.scala 83:21]
  reg [31:0] regs_4; // @[util.scala 83:21]
  reg [31:0] regs_5; // @[util.scala 83:21]
  reg [31:0] regs_6; // @[util.scala 83:21]
  reg [31:0] regs_7; // @[util.scala 83:21]
  reg [31:0] regs_8; // @[util.scala 83:21]
  reg [31:0] regs_9; // @[util.scala 83:21]
  reg [31:0] regs_10; // @[util.scala 83:21]
  reg [31:0] regs_11; // @[util.scala 83:21]
  reg [31:0] regs_12; // @[util.scala 83:21]
  reg [31:0] regs_13; // @[util.scala 83:21]
  reg [31:0] regs_14; // @[util.scala 83:21]
  reg [31:0] regs_15; // @[util.scala 83:21]
  reg [31:0] regs_16; // @[util.scala 83:21]
  reg [31:0] regs_17; // @[util.scala 83:21]
  reg [31:0] regs_18; // @[util.scala 83:21]
  reg [31:0] regs_19; // @[util.scala 83:21]
  reg [31:0] regs_20; // @[util.scala 83:21]
  reg [31:0] regs_21; // @[util.scala 83:21]
  reg [31:0] regs_22; // @[util.scala 83:21]
  reg [31:0] regs_23; // @[util.scala 83:21]
  reg [31:0] regs_24; // @[util.scala 83:21]
  reg [31:0] regs_25; // @[util.scala 83:21]
  reg [31:0] regs_26; // @[util.scala 83:21]
  reg [31:0] regs_27; // @[util.scala 83:21]
  reg [31:0] regs_28; // @[util.scala 83:21]
  reg [31:0] regs_29; // @[util.scala 83:21]
  reg [31:0] regs_30; // @[util.scala 83:21]
  reg [31:0] regs_31; // @[util.scala 83:21]
  wire [31:0] _GEN_1 = 5'h1 == io_rptr ? regs_1 : regs_0; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_2 = 5'h2 == io_rptr ? regs_2 : _GEN_1; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_3 = 5'h3 == io_rptr ? regs_3 : _GEN_2; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_4 = 5'h4 == io_rptr ? regs_4 : _GEN_3; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_5 = 5'h5 == io_rptr ? regs_5 : _GEN_4; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_6 = 5'h6 == io_rptr ? regs_6 : _GEN_5; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_7 = 5'h7 == io_rptr ? regs_7 : _GEN_6; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_8 = 5'h8 == io_rptr ? regs_8 : _GEN_7; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_9 = 5'h9 == io_rptr ? regs_9 : _GEN_8; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_10 = 5'ha == io_rptr ? regs_10 : _GEN_9; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_11 = 5'hb == io_rptr ? regs_11 : _GEN_10; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_12 = 5'hc == io_rptr ? regs_12 : _GEN_11; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_13 = 5'hd == io_rptr ? regs_13 : _GEN_12; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_14 = 5'he == io_rptr ? regs_14 : _GEN_13; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_15 = 5'hf == io_rptr ? regs_15 : _GEN_14; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_16 = 5'h10 == io_rptr ? regs_16 : _GEN_15; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_17 = 5'h11 == io_rptr ? regs_17 : _GEN_16; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_18 = 5'h12 == io_rptr ? regs_18 : _GEN_17; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_19 = 5'h13 == io_rptr ? regs_19 : _GEN_18; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_20 = 5'h14 == io_rptr ? regs_20 : _GEN_19; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_21 = 5'h15 == io_rptr ? regs_21 : _GEN_20; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_22 = 5'h16 == io_rptr ? regs_22 : _GEN_21; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_23 = 5'h17 == io_rptr ? regs_23 : _GEN_22; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_24 = 5'h18 == io_rptr ? regs_24 : _GEN_23; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_25 = 5'h19 == io_rptr ? regs_25 : _GEN_24; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_26 = 5'h1a == io_rptr ? regs_26 : _GEN_25; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_27 = 5'h1b == io_rptr ? regs_27 : _GEN_26; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_28 = 5'h1c == io_rptr ? regs_28 : _GEN_27; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_29 = 5'h1d == io_rptr ? regs_29 : _GEN_28; // @[util.scala 85:14 util.scala 85:14]
  wire [31:0] _GEN_30 = 5'h1e == io_rptr ? regs_30 : _GEN_29; // @[util.scala 85:14 util.scala 85:14]
  reg [4:0] counterValue; // @[Counter.scala 60:40]
  wire [4:0] _wrap_value_T_1 = counterValue + 5'h1; // @[Counter.scala 76:24]
  assign io_dataOut = 5'h1f == io_rptr ? regs_31 : _GEN_30; // @[util.scala 85:14 util.scala 85:14]
  assign io_wcount = counterValue; // @[util.scala 92:13]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 83:21]
      regs_0 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h0 == io_wptr) begin // @[util.scala 88:19]
        regs_0 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_1 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h1 == io_wptr) begin // @[util.scala 88:19]
        regs_1 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_2 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h2 == io_wptr) begin // @[util.scala 88:19]
        regs_2 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_3 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h3 == io_wptr) begin // @[util.scala 88:19]
        regs_3 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_4 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h4 == io_wptr) begin // @[util.scala 88:19]
        regs_4 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_5 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h5 == io_wptr) begin // @[util.scala 88:19]
        regs_5 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_6 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h6 == io_wptr) begin // @[util.scala 88:19]
        regs_6 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_7 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h7 == io_wptr) begin // @[util.scala 88:19]
        regs_7 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_8 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h8 == io_wptr) begin // @[util.scala 88:19]
        regs_8 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_9 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h9 == io_wptr) begin // @[util.scala 88:19]
        regs_9 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_10 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'ha == io_wptr) begin // @[util.scala 88:19]
        regs_10 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_11 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'hb == io_wptr) begin // @[util.scala 88:19]
        regs_11 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_12 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'hc == io_wptr) begin // @[util.scala 88:19]
        regs_12 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_13 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'hd == io_wptr) begin // @[util.scala 88:19]
        regs_13 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_14 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'he == io_wptr) begin // @[util.scala 88:19]
        regs_14 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_15 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'hf == io_wptr) begin // @[util.scala 88:19]
        regs_15 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_16 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h10 == io_wptr) begin // @[util.scala 88:19]
        regs_16 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_17 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h11 == io_wptr) begin // @[util.scala 88:19]
        regs_17 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_18 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h12 == io_wptr) begin // @[util.scala 88:19]
        regs_18 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_19 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h13 == io_wptr) begin // @[util.scala 88:19]
        regs_19 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_20 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h14 == io_wptr) begin // @[util.scala 88:19]
        regs_20 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_21 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h15 == io_wptr) begin // @[util.scala 88:19]
        regs_21 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_22 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h16 == io_wptr) begin // @[util.scala 88:19]
        regs_22 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_23 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h17 == io_wptr) begin // @[util.scala 88:19]
        regs_23 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_24 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h18 == io_wptr) begin // @[util.scala 88:19]
        regs_24 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_25 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h19 == io_wptr) begin // @[util.scala 88:19]
        regs_25 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_26 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h1a == io_wptr) begin // @[util.scala 88:19]
        regs_26 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_27 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h1b == io_wptr) begin // @[util.scala 88:19]
        regs_27 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_28 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h1c == io_wptr) begin // @[util.scala 88:19]
        regs_28 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_29 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h1d == io_wptr) begin // @[util.scala 88:19]
        regs_29 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_30 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h1e == io_wptr) begin // @[util.scala 88:19]
        regs_30 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[util.scala 83:21]
      regs_31 <= 32'h0; // @[util.scala 83:21]
    end else if (io_writeFlag) begin // @[util.scala 87:21]
      if (5'h1f == io_wptr) begin // @[util.scala 88:19]
        regs_31 <= io_dataIn; // @[util.scala 88:19]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      counterValue <= 5'h0; // @[Counter.scala 60:40]
    end else if (io_writeFlag) begin // @[Counter.scala 118:17]
      counterValue <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  counterValue = _RAND_32[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  input          io_start,
  input  [31:0]  io_root,
  output         io_issue_sync,
  input  [3:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 476:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 476:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 476:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 476:34]
  wire  edge_cache_clock; // @[BFS.scala 490:26]
  wire  edge_cache_reset; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 490:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 490:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 490:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 490:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 490:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 490:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 490:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 490:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 490:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 490:26]
  wire [4:0] edge_cache_io_free_ptr; // @[BFS.scala 490:26]
  wire [31:0] edge_cache_io_read_edge_num; // @[BFS.scala 490:26]
  wire  r_demux_aclk; // @[BFS.scala 493:23]
  wire  r_demux_aresetn; // @[BFS.scala 493:23]
  wire [127:0] r_demux_s_axis_tdata; // @[BFS.scala 493:23]
  wire [15:0] r_demux_s_axis_tkeep; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tlast; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tvalid; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tready; // @[BFS.scala 493:23]
  wire [5:0] r_demux_s_axis_tid; // @[BFS.scala 493:23]
  wire [255:0] r_demux_m_axis_tdata; // @[BFS.scala 493:23]
  wire [31:0] r_demux_m_axis_tkeep; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tlast; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tvalid; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tready; // @[BFS.scala 493:23]
  wire [11:0] r_demux_m_axis_tid; // @[BFS.scala 493:23]
  wire  arbi_clock; // @[BFS.scala 514:20]
  wire  arbi_reset; // @[BFS.scala 514:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 514:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 514:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 514:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 514:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 514:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 514:20]
  wire  arbi_io_out_ready; // @[BFS.scala 514:20]
  wire  arbi_io_out_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 514:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 514:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 514:20]
  wire  num_regfile_clock; // @[BFS.scala 528:27]
  wire  num_regfile_reset; // @[BFS.scala 528:27]
  wire [31:0] num_regfile_io_dataIn; // @[BFS.scala 528:27]
  wire [31:0] num_regfile_io_dataOut; // @[BFS.scala 528:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_wcount; // @[BFS.scala 528:27]
  wire  vertex_out_fifo_full; // @[BFS.scala 590:31]
  wire [131:0] vertex_out_fifo_din; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 590:31]
  wire [131:0] vertex_out_fifo_dout; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 590:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 590:31]
  reg [2:0] upward_status; // @[BFS.scala 469:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 470:30]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 471:35]
  wire [4:0] vertex_read_id_lo = vertex_read_buffer_data_count[4:0]; // @[BFS.scala 484:78 BFS.scala 484:78]
  wire  r_demux_out_0_valid = r_demux_m_axis_tvalid[0]; // @[BFS.scala 505:42]
  wire [5:0] r_demux_out_0_bits_rid = r_demux_m_axis_tid[5:0]; // @[BFS.scala 506:42]
  wire  r_demux_out_0_bits_rlast = r_demux_m_axis_tlast[0]; // @[BFS.scala 507:46]
  wire [127:0] r_demux_out_0_bits_rdata = r_demux_m_axis_tdata[127:0]; // @[BFS.scala 508:46]
  wire  r_demux_out_1_ready = edge_cache_io_in_ready; // @[BFS.scala 494:25 BFS.scala 512:20]
  wire  r_demux_out_0_ready = ~vertex_out_fifo_full; // @[BFS.scala 603:51]
  wire [37:0] _arbi_io_in_1_bits_araddr_T = {vertex_read_buffer_dout, 6'h0}; // @[BFS.scala 516:86]
  wire [63:0] _GEN_29 = {{26'd0}, _arbi_io_in_1_bits_araddr_T}; // @[BFS.scala 516:56]
  wire  _arbi_io_in_1_valid_T_3 = inflight_vtxs < 64'h20; // @[BFS.scala 517:116]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 523:96]
  reg [1:0] status; // @[BFS.scala 543:23]
  reg [31:0] num; // @[BFS.scala 544:20]
  wire  _T = status == 2'h0; // @[BFS.scala 545:15]
  wire  _T_4 = status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready; // @[BFS.scala 545:66]
  wire  _T_8 = status == 2'h2; // @[BFS.scala 553:22]
  wire  _T_9 = status == 2'h1; // @[BFS.scala 553:60]
  wire  _T_10 = status == 2'h2 | status == 2'h1; // @[BFS.scala 553:50]
  wire [31:0] _num_T_2 = num - 32'h4; // @[BFS.scala 569:18]
  wire [31:0] _num_T_6 = num > 32'h4 ? _num_T_2 : 32'h0; // @[BFS.scala 575:17]
  wire [31:0] _GEN_6 = r_demux_out_0_bits_rlast ? 32'h0 : _num_T_6; // @[BFS.scala 572:45 BFS.scala 573:11 BFS.scala 575:11]
  wire  _keep_0_T_3 = _T & r_demux_out_0_bits_rid[5]; // @[BFS.scala 582:33]
  wire  _keep_0_T_4 = num_regfile_io_dataOut > 32'h0; // @[BFS.scala 582:109]
  wire  _keep_0_T_6 = num > 32'h0; // @[BFS.scala 583:51]
  wire  _keep_0_T_10 = ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 584:36]
  wire  _keep_0_T_11 = _T & ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 584:33]
  wire [31:0] _keep_0_T_15 = r_demux_out_0_bits_rdata[63:32] + 32'h2; // @[BFS.scala 585:80]
  wire [2:0] _keep_0_T_22 = 3'h4 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_30 = {{29'd0}, _keep_0_T_22}; // @[BFS.scala 586:56]
  wire  _keep_0_T_23 = num > _GEN_30; // @[BFS.scala 586:56]
  wire  _keep_0_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_0_T_23; // @[Mux.scala 98:16]
  wire  _keep_0_T_26 = _T_8 ? _keep_0_T_6 : _keep_0_T_25; // @[Mux.scala 98:16]
  wire  keep_0 = _keep_0_T_3 ? _keep_0_T_4 : _keep_0_T_26; // @[Mux.scala 98:16]
  wire  _keep_1_T_4 = num_regfile_io_dataOut > 32'h1; // @[BFS.scala 582:109]
  wire  _keep_1_T_6 = num > 32'h1; // @[BFS.scala 583:51]
  wire [2:0] _keep_1_T_22 = 3'h5 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_31 = {{29'd0}, _keep_1_T_22}; // @[BFS.scala 586:56]
  wire  _keep_1_T_23 = num > _GEN_31; // @[BFS.scala 586:56]
  wire  _keep_1_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_1_T_23; // @[Mux.scala 98:16]
  wire  _keep_1_T_26 = _T_8 ? _keep_1_T_6 : _keep_1_T_25; // @[Mux.scala 98:16]
  wire  keep_1 = _keep_0_T_3 ? _keep_1_T_4 : _keep_1_T_26; // @[Mux.scala 98:16]
  wire  _keep_2_T_4 = num_regfile_io_dataOut > 32'h2; // @[BFS.scala 582:109]
  wire  _keep_2_T_6 = num > 32'h2; // @[BFS.scala 583:51]
  wire [2:0] _keep_2_T_22 = 3'h6 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_32 = {{29'd0}, _keep_2_T_22}; // @[BFS.scala 586:56]
  wire  _keep_2_T_23 = num > _GEN_32; // @[BFS.scala 586:56]
  wire  _keep_2_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_2_T_23; // @[Mux.scala 98:16]
  wire  _keep_2_T_26 = _T_8 ? _keep_2_T_6 : _keep_2_T_25; // @[Mux.scala 98:16]
  wire  keep_2 = _keep_0_T_3 ? _keep_2_T_4 : _keep_2_T_26; // @[Mux.scala 98:16]
  wire  _keep_3_T_4 = num_regfile_io_dataOut > 32'h3; // @[BFS.scala 582:109]
  wire  _keep_3_T_6 = num > 32'h3; // @[BFS.scala 583:51]
  wire  _keep_3_T_16 = _keep_0_T_15 > 32'h3; // @[BFS.scala 585:87]
  wire [2:0] _keep_3_T_22 = 3'h7 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_33 = {{29'd0}, _keep_3_T_22}; // @[BFS.scala 586:56]
  wire  _keep_3_T_23 = num > _GEN_33; // @[BFS.scala 586:56]
  wire  _keep_3_T_25 = _keep_0_T_11 ? _keep_3_T_16 : _T_9 & _keep_3_T_23; // @[Mux.scala 98:16]
  wire  _keep_3_T_26 = _T_8 ? _keep_3_T_6 : _keep_3_T_25; // @[Mux.scala 98:16]
  wire  keep_3 = _keep_0_T_3 ? _keep_3_T_4 : _keep_3_T_26; // @[Mux.scala 98:16]
  wire [131:0] _vertex_out_fifo_io_din_T = {r_demux_out_0_bits_rdata,keep_3,keep_2,keep_1,keep_0}; // @[Cat.scala 30:58]
  wire [35:0] _vertex_out_fifo_io_din_T_1 = {io_root,4'h1}; // @[Cat.scala 30:58]
  wire [131:0] _vertex_out_fifo_io_din_T_4 = _vertex_read_buffer_io_rd_en_T_2 ? 132'h800000001 :
    _vertex_out_fifo_io_din_T; // @[Mux.scala 98:16]
  reg  syncRecv_0; // @[BFS.scala 606:25]
  reg  syncRecv_1; // @[BFS.scala 606:25]
  reg  syncRecv_2; // @[BFS.scala 606:25]
  reg  syncRecv_3; // @[BFS.scala 606:25]
  wire  _GEN_10 = io_signal ? 1'h0 : syncRecv_0; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_11 = io_recv_sync[0] | _GEN_10; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_12 = io_signal ? 1'h0 : syncRecv_1; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_13 = io_recv_sync[1] | _GEN_12; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_14 = io_signal ? 1'h0 : syncRecv_2; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_15 = io_recv_sync[2] | _GEN_14; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_16 = io_signal ? 1'h0 : syncRecv_3; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_17 = io_recv_sync[3] | _GEN_16; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 616:34]
  wire [31:0] _T_46 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 112:12]
  wire  _T_50 = _T_46[0] & ~vertex_read_buffer_empty; // @[util.scala 112:36]
  wire [2:0] _GEN_19 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 629:53 BFS.scala 630:19 BFS.scala 469:30]
  wire [2:0] _GEN_20 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3) ? 3'h3 : _GEN_19; // @[BFS.scala 623:71]
  wire  _T_74 = r_demux_out_0_valid & r_demux_out_0_ready & _keep_0_T_10; // @[BFS.scala 635:77]
  wire [63:0] _GEN_35 = {{32'd0}, r_demux_out_0_bits_rdata[63:32]}; // @[BFS.scala 637:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_35; // @[BFS.scala 637:46]
  wire  _T_77 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 640:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 644:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 646:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 476:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 490:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_free_ptr(edge_cache_io_free_ptr),
    .io_read_edge_num(edge_cache_io_read_edge_num)
  );
  r_demux r_demux ( // @[BFS.scala 493:23]
    .aclk(r_demux_aclk),
    .aresetn(r_demux_aresetn),
    .s_axis_tdata(r_demux_s_axis_tdata),
    .s_axis_tkeep(r_demux_s_axis_tkeep),
    .s_axis_tlast(r_demux_s_axis_tlast),
    .s_axis_tvalid(r_demux_s_axis_tvalid),
    .s_axis_tready(r_demux_s_axis_tready),
    .s_axis_tid(r_demux_s_axis_tid),
    .m_axis_tdata(r_demux_m_axis_tdata),
    .m_axis_tkeep(r_demux_m_axis_tkeep),
    .m_axis_tlast(r_demux_m_axis_tlast),
    .m_axis_tvalid(r_demux_m_axis_tvalid),
    .m_axis_tready(r_demux_m_axis_tready),
    .m_axis_tid(r_demux_m_axis_tid)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 514:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  regFile num_regfile ( // @[BFS.scala 528:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr),
    .io_wcount(num_regfile_io_wcount)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 590:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 515:13]
  assign io_ddr_r_ready = r_demux_s_axis_tready; // @[BFS.scala 502:18]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 481:52]
  assign io_xbar_out_valid = vertex_out_fifo_valid; // @[BFS.scala 593:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_dout[131:4]; // @[BFS.scala 595:52]
  assign io_xbar_out_bits_tkeep = vertex_out_fifo_dout[3:0]; // @[BFS.scala 594:52]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 472:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 616:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 480:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 479:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 523:80]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 477:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 478:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = r_demux_m_axis_tvalid[1]; // @[BFS.scala 505:42]
  assign edge_cache_io_in_bits_rdata = r_demux_m_axis_tdata[255:128]; // @[BFS.scala 508:46]
  assign edge_cache_io_in_bits_rid = r_demux_m_axis_tid[11:6]; // @[BFS.scala 506:42]
  assign edge_cache_io_in_bits_rlast = r_demux_m_axis_tlast[1]; // @[BFS.scala 507:46]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 524:17]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 492:32]
  assign edge_cache_io_free_ptr = num_regfile_io_wcount; // @[BFS.scala 533:26]
  assign r_demux_aclk = clock; // @[BFS.scala 500:34]
  assign r_demux_aresetn = ~reset; // @[BFS.scala 501:25]
  assign r_demux_s_axis_tdata = io_ddr_r_bits_rdata; // @[BFS.scala 496:27]
  assign r_demux_s_axis_tkeep = 16'hffff; // @[nf_arm_doce_top.scala 117:85]
  assign r_demux_s_axis_tlast = io_ddr_r_bits_rlast; // @[BFS.scala 497:27]
  assign r_demux_s_axis_tvalid = io_ddr_r_valid; // @[BFS.scala 495:28]
  assign r_demux_s_axis_tid = io_ddr_r_bits_rid; // @[BFS.scala 499:25]
  assign r_demux_m_axis_tready = {r_demux_out_1_ready,r_demux_out_0_ready}; // @[BFS.scala 511:84]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 524:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & inflight_vtxs < 64'h20; // @[BFS.scala 517:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_29; // @[BFS.scala 516:56]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id_lo}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 515:13]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = edge_cache_io_read_edge_num; // @[BFS.scala 531:25]
  assign num_regfile_io_writeFlag = arbi_io_in_0_ready & arbi_io_in_0_valid; // @[BFS.scala 529:51]
  assign num_regfile_io_rptr = r_demux_out_0_bits_rid[4:0]; // @[BFS.scala 365:7]
  assign num_regfile_io_wptr = num_regfile_io_wcount; // @[BFS.scala 530:23]
  assign vertex_out_fifo_din = io_start ? {{96'd0}, _vertex_out_fifo_io_din_T_1} : _vertex_out_fifo_io_din_T_4; // @[Mux.scala 98:16]
  assign vertex_out_fifo_wr_en = r_demux_out_0_valid | _vertex_read_buffer_io_rd_en_T_2 | io_start; // @[BFS.scala 598:93]
  assign vertex_out_fifo_rd_en = io_xbar_out_ready; // @[BFS.scala 597:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 592:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 591:42]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 469:30]
      upward_status <= 3'h0; // @[BFS.scala 469:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 617:57]
      upward_status <= 3'h1; // @[BFS.scala 618:19]
    end else if (upward_status == 3'h1 & (_T_50 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3))) begin // @[BFS.scala 619:105]
      upward_status <= 3'h2; // @[BFS.scala 620:19]
    end else if (upward_status == 3'h2 & inflight_vtxs == 64'h0 & vertex_out_fifo_empty) begin // @[BFS.scala 621:110]
      upward_status <= 3'h4; // @[BFS.scala 622:19]
    end else begin
      upward_status <= _GEN_20;
    end
    if (reset) begin // @[BFS.scala 470:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 470:30]
    end else if (!(_T_77 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 641:91]
      if (_T_77) begin // @[BFS.scala 643:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 644:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 645:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 646:19]
      end
    end
    if (reset) begin // @[BFS.scala 471:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 471:35]
    end else if (io_signal) begin // @[BFS.scala 633:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 634:24]
    end else if (_T_74 & _T) begin // @[BFS.scala 636:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 637:24]
    end
    if (reset) begin // @[BFS.scala 543:23]
      status <= 2'h0; // @[BFS.scala 543:23]
    end else if (status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 545:99]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 546:45]
        status <= 2'h0; // @[BFS.scala 547:14]
      end else if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 548:61]
        status <= 2'h2; // @[BFS.scala 549:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 551:14]
      end
    end else if (_T_10 & r_demux_out_0_valid & r_demux_out_0_ready & r_demux_out_0_bits_rlast) begin // @[BFS.scala 554:117]
      status <= 2'h0; // @[BFS.scala 555:14]
    end
    if (reset) begin // @[BFS.scala 544:20]
      num <= 32'h0; // @[BFS.scala 544:20]
    end else if (_T_4 & ~r_demux_out_0_bits_rlast) begin // @[BFS.scala 559:112]
      if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 560:55]
        num <= num_regfile_io_dataOut; // @[BFS.scala 561:11]
      end else begin
        num <= r_demux_out_0_bits_rdata[63:32]; // @[BFS.scala 563:11]
      end
    end else if (_T_8 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 565:114]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 566:45]
        num <= 32'h0; // @[BFS.scala 567:11]
      end else begin
        num <= _num_T_2; // @[BFS.scala 569:11]
      end
    end else if (_T_9 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 571:119]
      num <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_0 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_1 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_2 <= _GEN_15;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_3 <= _GEN_17;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  status = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  num = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_3 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_1(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [3:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 476:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 476:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 476:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 476:34]
  wire  edge_cache_clock; // @[BFS.scala 490:26]
  wire  edge_cache_reset; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 490:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 490:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 490:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 490:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 490:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 490:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 490:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 490:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 490:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 490:26]
  wire [4:0] edge_cache_io_free_ptr; // @[BFS.scala 490:26]
  wire [31:0] edge_cache_io_read_edge_num; // @[BFS.scala 490:26]
  wire  r_demux_aclk; // @[BFS.scala 493:23]
  wire  r_demux_aresetn; // @[BFS.scala 493:23]
  wire [127:0] r_demux_s_axis_tdata; // @[BFS.scala 493:23]
  wire [15:0] r_demux_s_axis_tkeep; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tlast; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tvalid; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tready; // @[BFS.scala 493:23]
  wire [5:0] r_demux_s_axis_tid; // @[BFS.scala 493:23]
  wire [255:0] r_demux_m_axis_tdata; // @[BFS.scala 493:23]
  wire [31:0] r_demux_m_axis_tkeep; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tlast; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tvalid; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tready; // @[BFS.scala 493:23]
  wire [11:0] r_demux_m_axis_tid; // @[BFS.scala 493:23]
  wire  arbi_clock; // @[BFS.scala 514:20]
  wire  arbi_reset; // @[BFS.scala 514:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 514:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 514:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 514:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 514:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 514:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 514:20]
  wire  arbi_io_out_ready; // @[BFS.scala 514:20]
  wire  arbi_io_out_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 514:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 514:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 514:20]
  wire  num_regfile_clock; // @[BFS.scala 528:27]
  wire  num_regfile_reset; // @[BFS.scala 528:27]
  wire [31:0] num_regfile_io_dataIn; // @[BFS.scala 528:27]
  wire [31:0] num_regfile_io_dataOut; // @[BFS.scala 528:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_wcount; // @[BFS.scala 528:27]
  wire  vertex_out_fifo_full; // @[BFS.scala 590:31]
  wire [131:0] vertex_out_fifo_din; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 590:31]
  wire [131:0] vertex_out_fifo_dout; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 590:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 590:31]
  reg [2:0] upward_status; // @[BFS.scala 469:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 470:30]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 471:35]
  wire [4:0] vertex_read_id_lo = vertex_read_buffer_data_count[4:0]; // @[BFS.scala 484:78 BFS.scala 484:78]
  wire  r_demux_out_0_valid = r_demux_m_axis_tvalid[0]; // @[BFS.scala 505:42]
  wire [5:0] r_demux_out_0_bits_rid = r_demux_m_axis_tid[5:0]; // @[BFS.scala 506:42]
  wire  r_demux_out_0_bits_rlast = r_demux_m_axis_tlast[0]; // @[BFS.scala 507:46]
  wire [127:0] r_demux_out_0_bits_rdata = r_demux_m_axis_tdata[127:0]; // @[BFS.scala 508:46]
  wire  r_demux_out_1_ready = edge_cache_io_in_ready; // @[BFS.scala 494:25 BFS.scala 512:20]
  wire  r_demux_out_0_ready = ~vertex_out_fifo_full; // @[BFS.scala 603:51]
  wire [37:0] _arbi_io_in_1_bits_araddr_T = {vertex_read_buffer_dout, 6'h0}; // @[BFS.scala 516:86]
  wire [63:0] _GEN_29 = {{26'd0}, _arbi_io_in_1_bits_araddr_T}; // @[BFS.scala 516:56]
  wire  _arbi_io_in_1_valid_T_3 = inflight_vtxs < 64'h20; // @[BFS.scala 517:116]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 523:96]
  reg [1:0] status; // @[BFS.scala 543:23]
  reg [31:0] num; // @[BFS.scala 544:20]
  wire  _T = status == 2'h0; // @[BFS.scala 545:15]
  wire  _T_4 = status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready; // @[BFS.scala 545:66]
  wire  _T_8 = status == 2'h2; // @[BFS.scala 553:22]
  wire  _T_9 = status == 2'h1; // @[BFS.scala 553:60]
  wire  _T_10 = status == 2'h2 | status == 2'h1; // @[BFS.scala 553:50]
  wire [31:0] _num_T_2 = num - 32'h4; // @[BFS.scala 569:18]
  wire [31:0] _num_T_6 = num > 32'h4 ? _num_T_2 : 32'h0; // @[BFS.scala 575:17]
  wire [31:0] _GEN_6 = r_demux_out_0_bits_rlast ? 32'h0 : _num_T_6; // @[BFS.scala 572:45 BFS.scala 573:11 BFS.scala 575:11]
  wire  _keep_0_T_3 = _T & r_demux_out_0_bits_rid[5]; // @[BFS.scala 582:33]
  wire  _keep_0_T_4 = num_regfile_io_dataOut > 32'h0; // @[BFS.scala 582:109]
  wire  _keep_0_T_6 = num > 32'h0; // @[BFS.scala 583:51]
  wire  _keep_0_T_10 = ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 584:36]
  wire  _keep_0_T_11 = _T & ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 584:33]
  wire [31:0] _keep_0_T_15 = r_demux_out_0_bits_rdata[63:32] + 32'h2; // @[BFS.scala 585:80]
  wire [2:0] _keep_0_T_22 = 3'h4 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_30 = {{29'd0}, _keep_0_T_22}; // @[BFS.scala 586:56]
  wire  _keep_0_T_23 = num > _GEN_30; // @[BFS.scala 586:56]
  wire  _keep_0_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_0_T_23; // @[Mux.scala 98:16]
  wire  _keep_0_T_26 = _T_8 ? _keep_0_T_6 : _keep_0_T_25; // @[Mux.scala 98:16]
  wire  keep_0 = _keep_0_T_3 ? _keep_0_T_4 : _keep_0_T_26; // @[Mux.scala 98:16]
  wire  _keep_1_T_4 = num_regfile_io_dataOut > 32'h1; // @[BFS.scala 582:109]
  wire  _keep_1_T_6 = num > 32'h1; // @[BFS.scala 583:51]
  wire [2:0] _keep_1_T_22 = 3'h5 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_31 = {{29'd0}, _keep_1_T_22}; // @[BFS.scala 586:56]
  wire  _keep_1_T_23 = num > _GEN_31; // @[BFS.scala 586:56]
  wire  _keep_1_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_1_T_23; // @[Mux.scala 98:16]
  wire  _keep_1_T_26 = _T_8 ? _keep_1_T_6 : _keep_1_T_25; // @[Mux.scala 98:16]
  wire  keep_1 = _keep_0_T_3 ? _keep_1_T_4 : _keep_1_T_26; // @[Mux.scala 98:16]
  wire  _keep_2_T_4 = num_regfile_io_dataOut > 32'h2; // @[BFS.scala 582:109]
  wire  _keep_2_T_6 = num > 32'h2; // @[BFS.scala 583:51]
  wire [2:0] _keep_2_T_22 = 3'h6 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_32 = {{29'd0}, _keep_2_T_22}; // @[BFS.scala 586:56]
  wire  _keep_2_T_23 = num > _GEN_32; // @[BFS.scala 586:56]
  wire  _keep_2_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_2_T_23; // @[Mux.scala 98:16]
  wire  _keep_2_T_26 = _T_8 ? _keep_2_T_6 : _keep_2_T_25; // @[Mux.scala 98:16]
  wire  keep_2 = _keep_0_T_3 ? _keep_2_T_4 : _keep_2_T_26; // @[Mux.scala 98:16]
  wire  _keep_3_T_4 = num_regfile_io_dataOut > 32'h3; // @[BFS.scala 582:109]
  wire  _keep_3_T_6 = num > 32'h3; // @[BFS.scala 583:51]
  wire  _keep_3_T_16 = _keep_0_T_15 > 32'h3; // @[BFS.scala 585:87]
  wire [2:0] _keep_3_T_22 = 3'h7 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_33 = {{29'd0}, _keep_3_T_22}; // @[BFS.scala 586:56]
  wire  _keep_3_T_23 = num > _GEN_33; // @[BFS.scala 586:56]
  wire  _keep_3_T_25 = _keep_0_T_11 ? _keep_3_T_16 : _T_9 & _keep_3_T_23; // @[Mux.scala 98:16]
  wire  _keep_3_T_26 = _T_8 ? _keep_3_T_6 : _keep_3_T_25; // @[Mux.scala 98:16]
  wire  keep_3 = _keep_0_T_3 ? _keep_3_T_4 : _keep_3_T_26; // @[Mux.scala 98:16]
  wire [131:0] _vertex_out_fifo_io_din_T = {r_demux_out_0_bits_rdata,keep_3,keep_2,keep_1,keep_0}; // @[Cat.scala 30:58]
  reg  syncRecv_0; // @[BFS.scala 606:25]
  reg  syncRecv_1; // @[BFS.scala 606:25]
  reg  syncRecv_2; // @[BFS.scala 606:25]
  reg  syncRecv_3; // @[BFS.scala 606:25]
  wire  _GEN_10 = io_signal ? 1'h0 : syncRecv_0; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_11 = io_recv_sync[0] | _GEN_10; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_12 = io_signal ? 1'h0 : syncRecv_1; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_13 = io_recv_sync[1] | _GEN_12; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_14 = io_signal ? 1'h0 : syncRecv_2; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_15 = io_recv_sync[2] | _GEN_14; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_16 = io_signal ? 1'h0 : syncRecv_3; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_17 = io_recv_sync[3] | _GEN_16; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 616:34]
  wire [31:0] _T_46 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 112:12]
  wire  _T_50 = _T_46[0] & ~vertex_read_buffer_empty; // @[util.scala 112:36]
  wire [2:0] _GEN_19 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 629:53 BFS.scala 630:19 BFS.scala 469:30]
  wire [2:0] _GEN_20 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3) ? 3'h0 : _GEN_19; // @[BFS.scala 623:71]
  wire  _T_74 = r_demux_out_0_valid & r_demux_out_0_ready & _keep_0_T_10; // @[BFS.scala 635:77]
  wire [63:0] _GEN_35 = {{32'd0}, r_demux_out_0_bits_rdata[63:32]}; // @[BFS.scala 637:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_35; // @[BFS.scala 637:46]
  wire  _T_77 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 640:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 644:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 646:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 476:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 490:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_free_ptr(edge_cache_io_free_ptr),
    .io_read_edge_num(edge_cache_io_read_edge_num)
  );
  r_demux r_demux ( // @[BFS.scala 493:23]
    .aclk(r_demux_aclk),
    .aresetn(r_demux_aresetn),
    .s_axis_tdata(r_demux_s_axis_tdata),
    .s_axis_tkeep(r_demux_s_axis_tkeep),
    .s_axis_tlast(r_demux_s_axis_tlast),
    .s_axis_tvalid(r_demux_s_axis_tvalid),
    .s_axis_tready(r_demux_s_axis_tready),
    .s_axis_tid(r_demux_s_axis_tid),
    .m_axis_tdata(r_demux_m_axis_tdata),
    .m_axis_tkeep(r_demux_m_axis_tkeep),
    .m_axis_tlast(r_demux_m_axis_tlast),
    .m_axis_tvalid(r_demux_m_axis_tvalid),
    .m_axis_tready(r_demux_m_axis_tready),
    .m_axis_tid(r_demux_m_axis_tid)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 514:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  regFile num_regfile ( // @[BFS.scala 528:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr),
    .io_wcount(num_regfile_io_wcount)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 590:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 515:13]
  assign io_ddr_r_ready = r_demux_s_axis_tready; // @[BFS.scala 502:18]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 481:52]
  assign io_xbar_out_valid = vertex_out_fifo_valid; // @[BFS.scala 593:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_dout[131:4]; // @[BFS.scala 595:52]
  assign io_xbar_out_bits_tkeep = vertex_out_fifo_dout[3:0]; // @[BFS.scala 594:52]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 472:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 616:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 480:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 479:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 523:80]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 477:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 478:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = r_demux_m_axis_tvalid[1]; // @[BFS.scala 505:42]
  assign edge_cache_io_in_bits_rdata = r_demux_m_axis_tdata[255:128]; // @[BFS.scala 508:46]
  assign edge_cache_io_in_bits_rid = r_demux_m_axis_tid[11:6]; // @[BFS.scala 506:42]
  assign edge_cache_io_in_bits_rlast = r_demux_m_axis_tlast[1]; // @[BFS.scala 507:46]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 524:17]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 492:32]
  assign edge_cache_io_free_ptr = num_regfile_io_wcount; // @[BFS.scala 533:26]
  assign r_demux_aclk = clock; // @[BFS.scala 500:34]
  assign r_demux_aresetn = ~reset; // @[BFS.scala 501:25]
  assign r_demux_s_axis_tdata = io_ddr_r_bits_rdata; // @[BFS.scala 496:27]
  assign r_demux_s_axis_tkeep = 16'hffff; // @[nf_arm_doce_top.scala 117:85]
  assign r_demux_s_axis_tlast = io_ddr_r_bits_rlast; // @[BFS.scala 497:27]
  assign r_demux_s_axis_tvalid = io_ddr_r_valid; // @[BFS.scala 495:28]
  assign r_demux_s_axis_tid = io_ddr_r_bits_rid; // @[BFS.scala 499:25]
  assign r_demux_m_axis_tready = {r_demux_out_1_ready,r_demux_out_0_ready}; // @[BFS.scala 511:84]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 524:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & inflight_vtxs < 64'h20; // @[BFS.scala 517:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_29; // @[BFS.scala 516:56]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id_lo}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 515:13]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = edge_cache_io_read_edge_num; // @[BFS.scala 531:25]
  assign num_regfile_io_writeFlag = arbi_io_in_0_ready & arbi_io_in_0_valid; // @[BFS.scala 529:51]
  assign num_regfile_io_rptr = r_demux_out_0_bits_rid[4:0]; // @[BFS.scala 365:7]
  assign num_regfile_io_wptr = num_regfile_io_wcount; // @[BFS.scala 530:23]
  assign vertex_out_fifo_din = _vertex_read_buffer_io_rd_en_T_2 ? 132'h800000001 : _vertex_out_fifo_io_din_T; // @[Mux.scala 98:16]
  assign vertex_out_fifo_wr_en = r_demux_out_0_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 598:52]
  assign vertex_out_fifo_rd_en = io_xbar_out_ready; // @[BFS.scala 597:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 592:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 591:42]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 469:30]
      upward_status <= 3'h0; // @[BFS.scala 469:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 617:57]
      upward_status <= 3'h1; // @[BFS.scala 618:19]
    end else if (upward_status == 3'h1 & (_T_50 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3))) begin // @[BFS.scala 619:105]
      upward_status <= 3'h2; // @[BFS.scala 620:19]
    end else if (upward_status == 3'h2 & inflight_vtxs == 64'h0 & vertex_out_fifo_empty) begin // @[BFS.scala 621:110]
      upward_status <= 3'h4; // @[BFS.scala 622:19]
    end else begin
      upward_status <= _GEN_20;
    end
    if (reset) begin // @[BFS.scala 470:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 470:30]
    end else if (!(_T_77 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 641:91]
      if (_T_77) begin // @[BFS.scala 643:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 644:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 645:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 646:19]
      end
    end
    if (reset) begin // @[BFS.scala 471:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 471:35]
    end else if (io_signal) begin // @[BFS.scala 633:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 634:24]
    end else if (_T_74 & _T) begin // @[BFS.scala 636:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 637:24]
    end
    if (reset) begin // @[BFS.scala 543:23]
      status <= 2'h0; // @[BFS.scala 543:23]
    end else if (status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 545:99]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 546:45]
        status <= 2'h0; // @[BFS.scala 547:14]
      end else if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 548:61]
        status <= 2'h2; // @[BFS.scala 549:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 551:14]
      end
    end else if (_T_10 & r_demux_out_0_valid & r_demux_out_0_ready & r_demux_out_0_bits_rlast) begin // @[BFS.scala 554:117]
      status <= 2'h0; // @[BFS.scala 555:14]
    end
    if (reset) begin // @[BFS.scala 544:20]
      num <= 32'h0; // @[BFS.scala 544:20]
    end else if (_T_4 & ~r_demux_out_0_bits_rlast) begin // @[BFS.scala 559:112]
      if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 560:55]
        num <= num_regfile_io_dataOut; // @[BFS.scala 561:11]
      end else begin
        num <= r_demux_out_0_bits_rdata[63:32]; // @[BFS.scala 563:11]
      end
    end else if (_T_8 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 565:114]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 566:45]
        num <= 32'h0; // @[BFS.scala 567:11]
      end else begin
        num <= _num_T_2; // @[BFS.scala 569:11]
      end
    end else if (_T_9 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 571:119]
      num <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_0 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_1 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_2 <= _GEN_15;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_3 <= _GEN_17;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  status = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  num = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_3 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_2(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [3:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 476:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 476:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 476:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 476:34]
  wire  edge_cache_clock; // @[BFS.scala 490:26]
  wire  edge_cache_reset; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 490:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 490:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 490:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 490:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 490:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 490:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 490:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 490:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 490:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 490:26]
  wire [4:0] edge_cache_io_free_ptr; // @[BFS.scala 490:26]
  wire [31:0] edge_cache_io_read_edge_num; // @[BFS.scala 490:26]
  wire  r_demux_aclk; // @[BFS.scala 493:23]
  wire  r_demux_aresetn; // @[BFS.scala 493:23]
  wire [127:0] r_demux_s_axis_tdata; // @[BFS.scala 493:23]
  wire [15:0] r_demux_s_axis_tkeep; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tlast; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tvalid; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tready; // @[BFS.scala 493:23]
  wire [5:0] r_demux_s_axis_tid; // @[BFS.scala 493:23]
  wire [255:0] r_demux_m_axis_tdata; // @[BFS.scala 493:23]
  wire [31:0] r_demux_m_axis_tkeep; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tlast; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tvalid; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tready; // @[BFS.scala 493:23]
  wire [11:0] r_demux_m_axis_tid; // @[BFS.scala 493:23]
  wire  arbi_clock; // @[BFS.scala 514:20]
  wire  arbi_reset; // @[BFS.scala 514:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 514:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 514:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 514:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 514:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 514:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 514:20]
  wire  arbi_io_out_ready; // @[BFS.scala 514:20]
  wire  arbi_io_out_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 514:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 514:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 514:20]
  wire  num_regfile_clock; // @[BFS.scala 528:27]
  wire  num_regfile_reset; // @[BFS.scala 528:27]
  wire [31:0] num_regfile_io_dataIn; // @[BFS.scala 528:27]
  wire [31:0] num_regfile_io_dataOut; // @[BFS.scala 528:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_wcount; // @[BFS.scala 528:27]
  wire  vertex_out_fifo_full; // @[BFS.scala 590:31]
  wire [131:0] vertex_out_fifo_din; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 590:31]
  wire [131:0] vertex_out_fifo_dout; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 590:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 590:31]
  reg [2:0] upward_status; // @[BFS.scala 469:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 470:30]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 471:35]
  wire [4:0] vertex_read_id_lo = vertex_read_buffer_data_count[4:0]; // @[BFS.scala 484:78 BFS.scala 484:78]
  wire  r_demux_out_0_valid = r_demux_m_axis_tvalid[0]; // @[BFS.scala 505:42]
  wire [5:0] r_demux_out_0_bits_rid = r_demux_m_axis_tid[5:0]; // @[BFS.scala 506:42]
  wire  r_demux_out_0_bits_rlast = r_demux_m_axis_tlast[0]; // @[BFS.scala 507:46]
  wire [127:0] r_demux_out_0_bits_rdata = r_demux_m_axis_tdata[127:0]; // @[BFS.scala 508:46]
  wire  r_demux_out_1_ready = edge_cache_io_in_ready; // @[BFS.scala 494:25 BFS.scala 512:20]
  wire  r_demux_out_0_ready = ~vertex_out_fifo_full; // @[BFS.scala 603:51]
  wire [37:0] _arbi_io_in_1_bits_araddr_T = {vertex_read_buffer_dout, 6'h0}; // @[BFS.scala 516:86]
  wire [63:0] _GEN_29 = {{26'd0}, _arbi_io_in_1_bits_araddr_T}; // @[BFS.scala 516:56]
  wire  _arbi_io_in_1_valid_T_3 = inflight_vtxs < 64'h20; // @[BFS.scala 517:116]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 523:96]
  reg [1:0] status; // @[BFS.scala 543:23]
  reg [31:0] num; // @[BFS.scala 544:20]
  wire  _T = status == 2'h0; // @[BFS.scala 545:15]
  wire  _T_4 = status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready; // @[BFS.scala 545:66]
  wire  _T_8 = status == 2'h2; // @[BFS.scala 553:22]
  wire  _T_9 = status == 2'h1; // @[BFS.scala 553:60]
  wire  _T_10 = status == 2'h2 | status == 2'h1; // @[BFS.scala 553:50]
  wire [31:0] _num_T_2 = num - 32'h4; // @[BFS.scala 569:18]
  wire [31:0] _num_T_6 = num > 32'h4 ? _num_T_2 : 32'h0; // @[BFS.scala 575:17]
  wire [31:0] _GEN_6 = r_demux_out_0_bits_rlast ? 32'h0 : _num_T_6; // @[BFS.scala 572:45 BFS.scala 573:11 BFS.scala 575:11]
  wire  _keep_0_T_3 = _T & r_demux_out_0_bits_rid[5]; // @[BFS.scala 582:33]
  wire  _keep_0_T_4 = num_regfile_io_dataOut > 32'h0; // @[BFS.scala 582:109]
  wire  _keep_0_T_6 = num > 32'h0; // @[BFS.scala 583:51]
  wire  _keep_0_T_10 = ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 584:36]
  wire  _keep_0_T_11 = _T & ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 584:33]
  wire [31:0] _keep_0_T_15 = r_demux_out_0_bits_rdata[63:32] + 32'h2; // @[BFS.scala 585:80]
  wire [2:0] _keep_0_T_22 = 3'h4 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_30 = {{29'd0}, _keep_0_T_22}; // @[BFS.scala 586:56]
  wire  _keep_0_T_23 = num > _GEN_30; // @[BFS.scala 586:56]
  wire  _keep_0_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_0_T_23; // @[Mux.scala 98:16]
  wire  _keep_0_T_26 = _T_8 ? _keep_0_T_6 : _keep_0_T_25; // @[Mux.scala 98:16]
  wire  keep_0 = _keep_0_T_3 ? _keep_0_T_4 : _keep_0_T_26; // @[Mux.scala 98:16]
  wire  _keep_1_T_4 = num_regfile_io_dataOut > 32'h1; // @[BFS.scala 582:109]
  wire  _keep_1_T_6 = num > 32'h1; // @[BFS.scala 583:51]
  wire [2:0] _keep_1_T_22 = 3'h5 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_31 = {{29'd0}, _keep_1_T_22}; // @[BFS.scala 586:56]
  wire  _keep_1_T_23 = num > _GEN_31; // @[BFS.scala 586:56]
  wire  _keep_1_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_1_T_23; // @[Mux.scala 98:16]
  wire  _keep_1_T_26 = _T_8 ? _keep_1_T_6 : _keep_1_T_25; // @[Mux.scala 98:16]
  wire  keep_1 = _keep_0_T_3 ? _keep_1_T_4 : _keep_1_T_26; // @[Mux.scala 98:16]
  wire  _keep_2_T_4 = num_regfile_io_dataOut > 32'h2; // @[BFS.scala 582:109]
  wire  _keep_2_T_6 = num > 32'h2; // @[BFS.scala 583:51]
  wire [2:0] _keep_2_T_22 = 3'h6 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_32 = {{29'd0}, _keep_2_T_22}; // @[BFS.scala 586:56]
  wire  _keep_2_T_23 = num > _GEN_32; // @[BFS.scala 586:56]
  wire  _keep_2_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_2_T_23; // @[Mux.scala 98:16]
  wire  _keep_2_T_26 = _T_8 ? _keep_2_T_6 : _keep_2_T_25; // @[Mux.scala 98:16]
  wire  keep_2 = _keep_0_T_3 ? _keep_2_T_4 : _keep_2_T_26; // @[Mux.scala 98:16]
  wire  _keep_3_T_4 = num_regfile_io_dataOut > 32'h3; // @[BFS.scala 582:109]
  wire  _keep_3_T_6 = num > 32'h3; // @[BFS.scala 583:51]
  wire  _keep_3_T_16 = _keep_0_T_15 > 32'h3; // @[BFS.scala 585:87]
  wire [2:0] _keep_3_T_22 = 3'h7 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_33 = {{29'd0}, _keep_3_T_22}; // @[BFS.scala 586:56]
  wire  _keep_3_T_23 = num > _GEN_33; // @[BFS.scala 586:56]
  wire  _keep_3_T_25 = _keep_0_T_11 ? _keep_3_T_16 : _T_9 & _keep_3_T_23; // @[Mux.scala 98:16]
  wire  _keep_3_T_26 = _T_8 ? _keep_3_T_6 : _keep_3_T_25; // @[Mux.scala 98:16]
  wire  keep_3 = _keep_0_T_3 ? _keep_3_T_4 : _keep_3_T_26; // @[Mux.scala 98:16]
  wire [131:0] _vertex_out_fifo_io_din_T = {r_demux_out_0_bits_rdata,keep_3,keep_2,keep_1,keep_0}; // @[Cat.scala 30:58]
  reg  syncRecv_0; // @[BFS.scala 606:25]
  reg  syncRecv_1; // @[BFS.scala 606:25]
  reg  syncRecv_2; // @[BFS.scala 606:25]
  reg  syncRecv_3; // @[BFS.scala 606:25]
  wire  _GEN_10 = io_signal ? 1'h0 : syncRecv_0; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_11 = io_recv_sync[0] | _GEN_10; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_12 = io_signal ? 1'h0 : syncRecv_1; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_13 = io_recv_sync[1] | _GEN_12; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_14 = io_signal ? 1'h0 : syncRecv_2; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_15 = io_recv_sync[2] | _GEN_14; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_16 = io_signal ? 1'h0 : syncRecv_3; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_17 = io_recv_sync[3] | _GEN_16; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 616:34]
  wire [31:0] _T_46 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 112:12]
  wire  _T_50 = _T_46[0] & ~vertex_read_buffer_empty; // @[util.scala 112:36]
  wire [2:0] _GEN_19 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 629:53 BFS.scala 630:19 BFS.scala 469:30]
  wire [2:0] _GEN_20 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3) ? 3'h0 : _GEN_19; // @[BFS.scala 623:71]
  wire  _T_74 = r_demux_out_0_valid & r_demux_out_0_ready & _keep_0_T_10; // @[BFS.scala 635:77]
  wire [63:0] _GEN_35 = {{32'd0}, r_demux_out_0_bits_rdata[63:32]}; // @[BFS.scala 637:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_35; // @[BFS.scala 637:46]
  wire  _T_77 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 640:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 644:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 646:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 476:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 490:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_free_ptr(edge_cache_io_free_ptr),
    .io_read_edge_num(edge_cache_io_read_edge_num)
  );
  r_demux r_demux ( // @[BFS.scala 493:23]
    .aclk(r_demux_aclk),
    .aresetn(r_demux_aresetn),
    .s_axis_tdata(r_demux_s_axis_tdata),
    .s_axis_tkeep(r_demux_s_axis_tkeep),
    .s_axis_tlast(r_demux_s_axis_tlast),
    .s_axis_tvalid(r_demux_s_axis_tvalid),
    .s_axis_tready(r_demux_s_axis_tready),
    .s_axis_tid(r_demux_s_axis_tid),
    .m_axis_tdata(r_demux_m_axis_tdata),
    .m_axis_tkeep(r_demux_m_axis_tkeep),
    .m_axis_tlast(r_demux_m_axis_tlast),
    .m_axis_tvalid(r_demux_m_axis_tvalid),
    .m_axis_tready(r_demux_m_axis_tready),
    .m_axis_tid(r_demux_m_axis_tid)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 514:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  regFile num_regfile ( // @[BFS.scala 528:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr),
    .io_wcount(num_regfile_io_wcount)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 590:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 515:13]
  assign io_ddr_r_ready = r_demux_s_axis_tready; // @[BFS.scala 502:18]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 481:52]
  assign io_xbar_out_valid = vertex_out_fifo_valid; // @[BFS.scala 593:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_dout[131:4]; // @[BFS.scala 595:52]
  assign io_xbar_out_bits_tkeep = vertex_out_fifo_dout[3:0]; // @[BFS.scala 594:52]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 472:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 616:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 480:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 479:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 523:80]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 477:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 478:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = r_demux_m_axis_tvalid[1]; // @[BFS.scala 505:42]
  assign edge_cache_io_in_bits_rdata = r_demux_m_axis_tdata[255:128]; // @[BFS.scala 508:46]
  assign edge_cache_io_in_bits_rid = r_demux_m_axis_tid[11:6]; // @[BFS.scala 506:42]
  assign edge_cache_io_in_bits_rlast = r_demux_m_axis_tlast[1]; // @[BFS.scala 507:46]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 524:17]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 492:32]
  assign edge_cache_io_free_ptr = num_regfile_io_wcount; // @[BFS.scala 533:26]
  assign r_demux_aclk = clock; // @[BFS.scala 500:34]
  assign r_demux_aresetn = ~reset; // @[BFS.scala 501:25]
  assign r_demux_s_axis_tdata = io_ddr_r_bits_rdata; // @[BFS.scala 496:27]
  assign r_demux_s_axis_tkeep = 16'hffff; // @[nf_arm_doce_top.scala 117:85]
  assign r_demux_s_axis_tlast = io_ddr_r_bits_rlast; // @[BFS.scala 497:27]
  assign r_demux_s_axis_tvalid = io_ddr_r_valid; // @[BFS.scala 495:28]
  assign r_demux_s_axis_tid = io_ddr_r_bits_rid; // @[BFS.scala 499:25]
  assign r_demux_m_axis_tready = {r_demux_out_1_ready,r_demux_out_0_ready}; // @[BFS.scala 511:84]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 524:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & inflight_vtxs < 64'h20; // @[BFS.scala 517:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_29; // @[BFS.scala 516:56]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id_lo}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 515:13]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = edge_cache_io_read_edge_num; // @[BFS.scala 531:25]
  assign num_regfile_io_writeFlag = arbi_io_in_0_ready & arbi_io_in_0_valid; // @[BFS.scala 529:51]
  assign num_regfile_io_rptr = r_demux_out_0_bits_rid[4:0]; // @[BFS.scala 365:7]
  assign num_regfile_io_wptr = num_regfile_io_wcount; // @[BFS.scala 530:23]
  assign vertex_out_fifo_din = _vertex_read_buffer_io_rd_en_T_2 ? 132'h800000001 : _vertex_out_fifo_io_din_T; // @[Mux.scala 98:16]
  assign vertex_out_fifo_wr_en = r_demux_out_0_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 598:52]
  assign vertex_out_fifo_rd_en = io_xbar_out_ready; // @[BFS.scala 597:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 592:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 591:42]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 469:30]
      upward_status <= 3'h0; // @[BFS.scala 469:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 617:57]
      upward_status <= 3'h1; // @[BFS.scala 618:19]
    end else if (upward_status == 3'h1 & (_T_50 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3))) begin // @[BFS.scala 619:105]
      upward_status <= 3'h2; // @[BFS.scala 620:19]
    end else if (upward_status == 3'h2 & inflight_vtxs == 64'h0 & vertex_out_fifo_empty) begin // @[BFS.scala 621:110]
      upward_status <= 3'h4; // @[BFS.scala 622:19]
    end else begin
      upward_status <= _GEN_20;
    end
    if (reset) begin // @[BFS.scala 470:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 470:30]
    end else if (!(_T_77 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 641:91]
      if (_T_77) begin // @[BFS.scala 643:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 644:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 645:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 646:19]
      end
    end
    if (reset) begin // @[BFS.scala 471:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 471:35]
    end else if (io_signal) begin // @[BFS.scala 633:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 634:24]
    end else if (_T_74 & _T) begin // @[BFS.scala 636:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 637:24]
    end
    if (reset) begin // @[BFS.scala 543:23]
      status <= 2'h0; // @[BFS.scala 543:23]
    end else if (status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 545:99]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 546:45]
        status <= 2'h0; // @[BFS.scala 547:14]
      end else if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 548:61]
        status <= 2'h2; // @[BFS.scala 549:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 551:14]
      end
    end else if (_T_10 & r_demux_out_0_valid & r_demux_out_0_ready & r_demux_out_0_bits_rlast) begin // @[BFS.scala 554:117]
      status <= 2'h0; // @[BFS.scala 555:14]
    end
    if (reset) begin // @[BFS.scala 544:20]
      num <= 32'h0; // @[BFS.scala 544:20]
    end else if (_T_4 & ~r_demux_out_0_bits_rlast) begin // @[BFS.scala 559:112]
      if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 560:55]
        num <= num_regfile_io_dataOut; // @[BFS.scala 561:11]
      end else begin
        num <= r_demux_out_0_bits_rdata[63:32]; // @[BFS.scala 563:11]
      end
    end else if (_T_8 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 565:114]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 566:45]
        num <= 32'h0; // @[BFS.scala 567:11]
      end else begin
        num <= _num_T_2; // @[BFS.scala 569:11]
      end
    end else if (_T_9 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 571:119]
      num <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_0 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_1 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_2 <= _GEN_15;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_3 <= _GEN_17;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  status = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  num = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_3 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_3(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [3:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 476:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 476:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 476:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 476:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 476:34]
  wire  edge_cache_clock; // @[BFS.scala 490:26]
  wire  edge_cache_reset; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 490:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 490:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 490:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 490:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 490:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 490:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 490:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 490:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 490:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 490:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 490:26]
  wire [4:0] edge_cache_io_free_ptr; // @[BFS.scala 490:26]
  wire [31:0] edge_cache_io_read_edge_num; // @[BFS.scala 490:26]
  wire  r_demux_aclk; // @[BFS.scala 493:23]
  wire  r_demux_aresetn; // @[BFS.scala 493:23]
  wire [127:0] r_demux_s_axis_tdata; // @[BFS.scala 493:23]
  wire [15:0] r_demux_s_axis_tkeep; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tlast; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tvalid; // @[BFS.scala 493:23]
  wire  r_demux_s_axis_tready; // @[BFS.scala 493:23]
  wire [5:0] r_demux_s_axis_tid; // @[BFS.scala 493:23]
  wire [255:0] r_demux_m_axis_tdata; // @[BFS.scala 493:23]
  wire [31:0] r_demux_m_axis_tkeep; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tlast; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tvalid; // @[BFS.scala 493:23]
  wire [1:0] r_demux_m_axis_tready; // @[BFS.scala 493:23]
  wire [11:0] r_demux_m_axis_tid; // @[BFS.scala 493:23]
  wire  arbi_clock; // @[BFS.scala 514:20]
  wire  arbi_reset; // @[BFS.scala 514:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 514:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 514:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 514:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 514:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 514:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 514:20]
  wire  arbi_io_out_ready; // @[BFS.scala 514:20]
  wire  arbi_io_out_valid; // @[BFS.scala 514:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 514:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 514:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 514:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 514:20]
  wire  num_regfile_clock; // @[BFS.scala 528:27]
  wire  num_regfile_reset; // @[BFS.scala 528:27]
  wire [31:0] num_regfile_io_dataIn; // @[BFS.scala 528:27]
  wire [31:0] num_regfile_io_dataOut; // @[BFS.scala 528:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 528:27]
  wire [4:0] num_regfile_io_wcount; // @[BFS.scala 528:27]
  wire  vertex_out_fifo_full; // @[BFS.scala 590:31]
  wire [131:0] vertex_out_fifo_din; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 590:31]
  wire [131:0] vertex_out_fifo_dout; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 590:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 590:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 590:31]
  reg [2:0] upward_status; // @[BFS.scala 469:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 470:30]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 471:35]
  wire [4:0] vertex_read_id_lo = vertex_read_buffer_data_count[4:0]; // @[BFS.scala 484:78 BFS.scala 484:78]
  wire  r_demux_out_0_valid = r_demux_m_axis_tvalid[0]; // @[BFS.scala 505:42]
  wire [5:0] r_demux_out_0_bits_rid = r_demux_m_axis_tid[5:0]; // @[BFS.scala 506:42]
  wire  r_demux_out_0_bits_rlast = r_demux_m_axis_tlast[0]; // @[BFS.scala 507:46]
  wire [127:0] r_demux_out_0_bits_rdata = r_demux_m_axis_tdata[127:0]; // @[BFS.scala 508:46]
  wire  r_demux_out_1_ready = edge_cache_io_in_ready; // @[BFS.scala 494:25 BFS.scala 512:20]
  wire  r_demux_out_0_ready = ~vertex_out_fifo_full; // @[BFS.scala 603:51]
  wire [37:0] _arbi_io_in_1_bits_araddr_T = {vertex_read_buffer_dout, 6'h0}; // @[BFS.scala 516:86]
  wire [63:0] _GEN_29 = {{26'd0}, _arbi_io_in_1_bits_araddr_T}; // @[BFS.scala 516:56]
  wire  _arbi_io_in_1_valid_T_3 = inflight_vtxs < 64'h20; // @[BFS.scala 517:116]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 523:96]
  reg [1:0] status; // @[BFS.scala 543:23]
  reg [31:0] num; // @[BFS.scala 544:20]
  wire  _T = status == 2'h0; // @[BFS.scala 545:15]
  wire  _T_4 = status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready; // @[BFS.scala 545:66]
  wire  _T_8 = status == 2'h2; // @[BFS.scala 553:22]
  wire  _T_9 = status == 2'h1; // @[BFS.scala 553:60]
  wire  _T_10 = status == 2'h2 | status == 2'h1; // @[BFS.scala 553:50]
  wire [31:0] _num_T_2 = num - 32'h4; // @[BFS.scala 569:18]
  wire [31:0] _num_T_6 = num > 32'h4 ? _num_T_2 : 32'h0; // @[BFS.scala 575:17]
  wire [31:0] _GEN_6 = r_demux_out_0_bits_rlast ? 32'h0 : _num_T_6; // @[BFS.scala 572:45 BFS.scala 573:11 BFS.scala 575:11]
  wire  _keep_0_T_3 = _T & r_demux_out_0_bits_rid[5]; // @[BFS.scala 582:33]
  wire  _keep_0_T_4 = num_regfile_io_dataOut > 32'h0; // @[BFS.scala 582:109]
  wire  _keep_0_T_6 = num > 32'h0; // @[BFS.scala 583:51]
  wire  _keep_0_T_10 = ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 584:36]
  wire  _keep_0_T_11 = _T & ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 584:33]
  wire [31:0] _keep_0_T_15 = r_demux_out_0_bits_rdata[63:32] + 32'h2; // @[BFS.scala 585:80]
  wire [2:0] _keep_0_T_22 = 3'h4 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_30 = {{29'd0}, _keep_0_T_22}; // @[BFS.scala 586:56]
  wire  _keep_0_T_23 = num > _GEN_30; // @[BFS.scala 586:56]
  wire  _keep_0_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_0_T_23; // @[Mux.scala 98:16]
  wire  _keep_0_T_26 = _T_8 ? _keep_0_T_6 : _keep_0_T_25; // @[Mux.scala 98:16]
  wire  keep_0 = _keep_0_T_3 ? _keep_0_T_4 : _keep_0_T_26; // @[Mux.scala 98:16]
  wire  _keep_1_T_4 = num_regfile_io_dataOut > 32'h1; // @[BFS.scala 582:109]
  wire  _keep_1_T_6 = num > 32'h1; // @[BFS.scala 583:51]
  wire [2:0] _keep_1_T_22 = 3'h5 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_31 = {{29'd0}, _keep_1_T_22}; // @[BFS.scala 586:56]
  wire  _keep_1_T_23 = num > _GEN_31; // @[BFS.scala 586:56]
  wire  _keep_1_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_1_T_23; // @[Mux.scala 98:16]
  wire  _keep_1_T_26 = _T_8 ? _keep_1_T_6 : _keep_1_T_25; // @[Mux.scala 98:16]
  wire  keep_1 = _keep_0_T_3 ? _keep_1_T_4 : _keep_1_T_26; // @[Mux.scala 98:16]
  wire  _keep_2_T_4 = num_regfile_io_dataOut > 32'h2; // @[BFS.scala 582:109]
  wire  _keep_2_T_6 = num > 32'h2; // @[BFS.scala 583:51]
  wire [2:0] _keep_2_T_22 = 3'h6 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_32 = {{29'd0}, _keep_2_T_22}; // @[BFS.scala 586:56]
  wire  _keep_2_T_23 = num > _GEN_32; // @[BFS.scala 586:56]
  wire  _keep_2_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_2_T_23; // @[Mux.scala 98:16]
  wire  _keep_2_T_26 = _T_8 ? _keep_2_T_6 : _keep_2_T_25; // @[Mux.scala 98:16]
  wire  keep_2 = _keep_0_T_3 ? _keep_2_T_4 : _keep_2_T_26; // @[Mux.scala 98:16]
  wire  _keep_3_T_4 = num_regfile_io_dataOut > 32'h3; // @[BFS.scala 582:109]
  wire  _keep_3_T_6 = num > 32'h3; // @[BFS.scala 583:51]
  wire  _keep_3_T_16 = _keep_0_T_15 > 32'h3; // @[BFS.scala 585:87]
  wire [2:0] _keep_3_T_22 = 3'h7 - 3'h2; // @[BFS.scala 586:78]
  wire [31:0] _GEN_33 = {{29'd0}, _keep_3_T_22}; // @[BFS.scala 586:56]
  wire  _keep_3_T_23 = num > _GEN_33; // @[BFS.scala 586:56]
  wire  _keep_3_T_25 = _keep_0_T_11 ? _keep_3_T_16 : _T_9 & _keep_3_T_23; // @[Mux.scala 98:16]
  wire  _keep_3_T_26 = _T_8 ? _keep_3_T_6 : _keep_3_T_25; // @[Mux.scala 98:16]
  wire  keep_3 = _keep_0_T_3 ? _keep_3_T_4 : _keep_3_T_26; // @[Mux.scala 98:16]
  wire [131:0] _vertex_out_fifo_io_din_T = {r_demux_out_0_bits_rdata,keep_3,keep_2,keep_1,keep_0}; // @[Cat.scala 30:58]
  reg  syncRecv_0; // @[BFS.scala 606:25]
  reg  syncRecv_1; // @[BFS.scala 606:25]
  reg  syncRecv_2; // @[BFS.scala 606:25]
  reg  syncRecv_3; // @[BFS.scala 606:25]
  wire  _GEN_10 = io_signal ? 1'h0 : syncRecv_0; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_11 = io_recv_sync[0] | _GEN_10; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_12 = io_signal ? 1'h0 : syncRecv_1; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_13 = io_recv_sync[1] | _GEN_12; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_14 = io_signal ? 1'h0 : syncRecv_2; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_15 = io_recv_sync[2] | _GEN_14; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _GEN_16 = io_signal ? 1'h0 : syncRecv_3; // @[BFS.scala 611:28 BFS.scala 612:11 BFS.scala 606:25]
  wire  _GEN_17 = io_recv_sync[3] | _GEN_16; // @[BFS.scala 609:28 BFS.scala 610:11]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 616:34]
  wire [31:0] _T_46 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 112:12]
  wire  _T_50 = _T_46[0] & ~vertex_read_buffer_empty; // @[util.scala 112:36]
  wire [2:0] _GEN_19 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 629:53 BFS.scala 630:19 BFS.scala 469:30]
  wire [2:0] _GEN_20 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3) ? 3'h0 : _GEN_19; // @[BFS.scala 623:71]
  wire  _T_74 = r_demux_out_0_valid & r_demux_out_0_ready & _keep_0_T_10; // @[BFS.scala 635:77]
  wire [63:0] _GEN_35 = {{32'd0}, r_demux_out_0_bits_rdata[63:32]}; // @[BFS.scala 637:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_35; // @[BFS.scala 637:46]
  wire  _T_77 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 640:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 644:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 646:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 476:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 490:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_free_ptr(edge_cache_io_free_ptr),
    .io_read_edge_num(edge_cache_io_read_edge_num)
  );
  r_demux r_demux ( // @[BFS.scala 493:23]
    .aclk(r_demux_aclk),
    .aresetn(r_demux_aresetn),
    .s_axis_tdata(r_demux_s_axis_tdata),
    .s_axis_tkeep(r_demux_s_axis_tkeep),
    .s_axis_tlast(r_demux_s_axis_tlast),
    .s_axis_tvalid(r_demux_s_axis_tvalid),
    .s_axis_tready(r_demux_s_axis_tready),
    .s_axis_tid(r_demux_s_axis_tid),
    .m_axis_tdata(r_demux_m_axis_tdata),
    .m_axis_tkeep(r_demux_m_axis_tkeep),
    .m_axis_tlast(r_demux_m_axis_tlast),
    .m_axis_tvalid(r_demux_m_axis_tvalid),
    .m_axis_tready(r_demux_m_axis_tready),
    .m_axis_tid(r_demux_m_axis_tid)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 514:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  regFile num_regfile ( // @[BFS.scala 528:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr),
    .io_wcount(num_regfile_io_wcount)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 590:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 515:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 515:13]
  assign io_ddr_r_ready = r_demux_s_axis_tready; // @[BFS.scala 502:18]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 481:52]
  assign io_xbar_out_valid = vertex_out_fifo_valid; // @[BFS.scala 593:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_dout[131:4]; // @[BFS.scala 595:52]
  assign io_xbar_out_bits_tkeep = vertex_out_fifo_dout[3:0]; // @[BFS.scala 594:52]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 472:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 616:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 480:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 479:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 523:80]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 477:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 478:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = r_demux_m_axis_tvalid[1]; // @[BFS.scala 505:42]
  assign edge_cache_io_in_bits_rdata = r_demux_m_axis_tdata[255:128]; // @[BFS.scala 508:46]
  assign edge_cache_io_in_bits_rid = r_demux_m_axis_tid[11:6]; // @[BFS.scala 506:42]
  assign edge_cache_io_in_bits_rlast = r_demux_m_axis_tlast[1]; // @[BFS.scala 507:46]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 524:17]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 492:32]
  assign edge_cache_io_free_ptr = num_regfile_io_wcount; // @[BFS.scala 533:26]
  assign r_demux_aclk = clock; // @[BFS.scala 500:34]
  assign r_demux_aresetn = ~reset; // @[BFS.scala 501:25]
  assign r_demux_s_axis_tdata = io_ddr_r_bits_rdata; // @[BFS.scala 496:27]
  assign r_demux_s_axis_tkeep = 16'hffff; // @[nf_arm_doce_top.scala 117:85]
  assign r_demux_s_axis_tlast = io_ddr_r_bits_rlast; // @[BFS.scala 497:27]
  assign r_demux_s_axis_tvalid = io_ddr_r_valid; // @[BFS.scala 495:28]
  assign r_demux_s_axis_tid = io_ddr_r_bits_rid; // @[BFS.scala 499:25]
  assign r_demux_m_axis_tready = {r_demux_out_1_ready,r_demux_out_0_ready}; // @[BFS.scala 511:84]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 524:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 524:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & inflight_vtxs < 64'h20; // @[BFS.scala 517:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_29; // @[BFS.scala 516:56]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id_lo}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 515:13]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = edge_cache_io_read_edge_num; // @[BFS.scala 531:25]
  assign num_regfile_io_writeFlag = arbi_io_in_0_ready & arbi_io_in_0_valid; // @[BFS.scala 529:51]
  assign num_regfile_io_rptr = r_demux_out_0_bits_rid[4:0]; // @[BFS.scala 365:7]
  assign num_regfile_io_wptr = num_regfile_io_wcount; // @[BFS.scala 530:23]
  assign vertex_out_fifo_din = _vertex_read_buffer_io_rd_en_T_2 ? 132'h800000001 : _vertex_out_fifo_io_din_T; // @[Mux.scala 98:16]
  assign vertex_out_fifo_wr_en = r_demux_out_0_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 598:52]
  assign vertex_out_fifo_rd_en = io_xbar_out_ready; // @[BFS.scala 597:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 592:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 591:42]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 469:30]
      upward_status <= 3'h0; // @[BFS.scala 469:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 617:57]
      upward_status <= 3'h1; // @[BFS.scala 618:19]
    end else if (upward_status == 3'h1 & (_T_50 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3))) begin // @[BFS.scala 619:105]
      upward_status <= 3'h2; // @[BFS.scala 620:19]
    end else if (upward_status == 3'h2 & inflight_vtxs == 64'h0 & vertex_out_fifo_empty) begin // @[BFS.scala 621:110]
      upward_status <= 3'h4; // @[BFS.scala 622:19]
    end else begin
      upward_status <= _GEN_20;
    end
    if (reset) begin // @[BFS.scala 470:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 470:30]
    end else if (!(_T_77 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 641:91]
      if (_T_77) begin // @[BFS.scala 643:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 644:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 645:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 646:19]
      end
    end
    if (reset) begin // @[BFS.scala 471:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 471:35]
    end else if (io_signal) begin // @[BFS.scala 633:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 634:24]
    end else if (_T_74 & _T) begin // @[BFS.scala 636:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 637:24]
    end
    if (reset) begin // @[BFS.scala 543:23]
      status <= 2'h0; // @[BFS.scala 543:23]
    end else if (status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 545:99]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 546:45]
        status <= 2'h0; // @[BFS.scala 547:14]
      end else if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 548:61]
        status <= 2'h2; // @[BFS.scala 549:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 551:14]
      end
    end else if (_T_10 & r_demux_out_0_valid & r_demux_out_0_ready & r_demux_out_0_bits_rlast) begin // @[BFS.scala 554:117]
      status <= 2'h0; // @[BFS.scala 555:14]
    end
    if (reset) begin // @[BFS.scala 544:20]
      num <= 32'h0; // @[BFS.scala 544:20]
    end else if (_T_4 & ~r_demux_out_0_bits_rlast) begin // @[BFS.scala 559:112]
      if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 560:55]
        num <= num_regfile_io_dataOut; // @[BFS.scala 561:11]
      end else begin
        num <= r_demux_out_0_bits_rdata[63:32]; // @[BFS.scala 563:11]
      end
    end else if (_T_8 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 565:114]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 566:45]
        num <= 32'h0; // @[BFS.scala 567:11]
      end else begin
        num <= _num_T_2; // @[BFS.scala 569:11]
      end
    end else if (_T_9 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 571:119]
      num <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_0 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_1 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_2 <= _GEN_15;
    end
    if (reset) begin // @[BFS.scala 606:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 606:25]
    end else begin
      syncRecv_3 <= _GEN_17;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  status = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  num = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_3 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module broadcast_xbar(
  input          clock,
  input          reset,
  output         io_ddr_in_0_ready,
  input          io_ddr_in_0_valid,
  input  [127:0] io_ddr_in_0_bits_tdata,
  input  [3:0]   io_ddr_in_0_bits_tkeep,
  output         io_ddr_in_1_ready,
  input          io_ddr_in_1_valid,
  input  [127:0] io_ddr_in_1_bits_tdata,
  input  [3:0]   io_ddr_in_1_bits_tkeep,
  output         io_ddr_in_2_ready,
  input          io_ddr_in_2_valid,
  input  [127:0] io_ddr_in_2_bits_tdata,
  input  [3:0]   io_ddr_in_2_bits_tkeep,
  output         io_ddr_in_3_ready,
  input          io_ddr_in_3_valid,
  input  [127:0] io_ddr_in_3_bits_tdata,
  input  [3:0]   io_ddr_in_3_bits_tkeep,
  input          io_pe_out_0_ready,
  output         io_pe_out_0_valid,
  output [511:0] io_pe_out_0_bits_tdata,
  output [15:0]  io_pe_out_0_bits_tkeep,
  input          io_pe_out_1_ready,
  output         io_pe_out_1_valid,
  output [511:0] io_pe_out_1_bits_tdata,
  output [15:0]  io_pe_out_1_bits_tkeep,
  input          io_pe_out_2_ready,
  output         io_pe_out_2_valid,
  output [511:0] io_pe_out_2_bits_tdata,
  output [15:0]  io_pe_out_2_bits_tkeep,
  input          io_pe_out_3_ready,
  output         io_pe_out_3_valid,
  output [511:0] io_pe_out_3_bits_tdata,
  output [15:0]  io_pe_out_3_bits_tkeep,
  input          io_pe_out_4_ready,
  output         io_pe_out_4_valid,
  output [511:0] io_pe_out_4_bits_tdata,
  output [15:0]  io_pe_out_4_bits_tkeep,
  input          io_pe_out_5_ready,
  output         io_pe_out_5_valid,
  output [511:0] io_pe_out_5_bits_tdata,
  output [15:0]  io_pe_out_5_bits_tkeep,
  input          io_pe_out_6_ready,
  output         io_pe_out_6_valid,
  output [511:0] io_pe_out_6_bits_tdata,
  output [15:0]  io_pe_out_6_bits_tkeep,
  input          io_pe_out_7_ready,
  output         io_pe_out_7_valid,
  output [511:0] io_pe_out_7_bits_tdata,
  output [15:0]  io_pe_out_7_bits_tkeep,
  input          io_pe_out_8_ready,
  output         io_pe_out_8_valid,
  output [511:0] io_pe_out_8_bits_tdata,
  output [15:0]  io_pe_out_8_bits_tkeep,
  input          io_pe_out_9_ready,
  output         io_pe_out_9_valid,
  output [511:0] io_pe_out_9_bits_tdata,
  output [15:0]  io_pe_out_9_bits_tkeep,
  input          io_pe_out_10_ready,
  output         io_pe_out_10_valid,
  output [511:0] io_pe_out_10_bits_tdata,
  output [15:0]  io_pe_out_10_bits_tkeep,
  input          io_pe_out_11_ready,
  output         io_pe_out_11_valid,
  output [511:0] io_pe_out_11_bits_tdata,
  output [15:0]  io_pe_out_11_bits_tkeep,
  input          io_pe_out_12_ready,
  output         io_pe_out_12_valid,
  output [511:0] io_pe_out_12_bits_tdata,
  output [15:0]  io_pe_out_12_bits_tkeep,
  input          io_pe_out_13_ready,
  output         io_pe_out_13_valid,
  output [511:0] io_pe_out_13_bits_tdata,
  output [15:0]  io_pe_out_13_bits_tkeep,
  input          io_pe_out_14_ready,
  output         io_pe_out_14_valid,
  output [511:0] io_pe_out_14_bits_tdata,
  output [15:0]  io_pe_out_14_bits_tkeep,
  input          io_pe_out_15_ready,
  output         io_pe_out_15_valid,
  output [511:0] io_pe_out_15_bits_tdata,
  output [15:0]  io_pe_out_15_bits_tkeep
);
  wire  xbar_aclk; // @[BFS.scala 660:20]
  wire  xbar_aresetn; // @[BFS.scala 660:20]
  wire [511:0] xbar_s_axis_tdata; // @[BFS.scala 660:20]
  wire [63:0] xbar_s_axis_tkeep; // @[BFS.scala 660:20]
  wire  xbar_s_axis_tlast; // @[BFS.scala 660:20]
  wire  xbar_s_axis_tvalid; // @[BFS.scala 660:20]
  wire  xbar_s_axis_tready; // @[BFS.scala 660:20]
  wire  xbar_s_axis_tid; // @[BFS.scala 660:20]
  wire [8191:0] xbar_m_axis_tdata; // @[BFS.scala 660:20]
  wire [1023:0] xbar_m_axis_tkeep; // @[BFS.scala 660:20]
  wire [15:0] xbar_m_axis_tlast; // @[BFS.scala 660:20]
  wire [15:0] xbar_m_axis_tvalid; // @[BFS.scala 660:20]
  wire [15:0] xbar_m_axis_tready; // @[BFS.scala 660:20]
  wire [15:0] xbar_m_axis_tid; // @[BFS.scala 660:20]
  wire  combiner_aclk; // @[BFS.scala 666:26]
  wire  combiner_aresetn; // @[BFS.scala 666:26]
  wire [511:0] combiner_s_axis_tdata; // @[BFS.scala 666:26]
  wire [63:0] combiner_s_axis_tkeep; // @[BFS.scala 666:26]
  wire [3:0] combiner_s_axis_tlast; // @[BFS.scala 666:26]
  wire [3:0] combiner_s_axis_tvalid; // @[BFS.scala 666:26]
  wire [3:0] combiner_s_axis_tready; // @[BFS.scala 666:26]
  wire [3:0] combiner_s_axis_tid; // @[BFS.scala 666:26]
  wire [511:0] combiner_m_axis_tdata; // @[BFS.scala 666:26]
  wire [63:0] combiner_m_axis_tkeep; // @[BFS.scala 666:26]
  wire  combiner_m_axis_tlast; // @[BFS.scala 666:26]
  wire  combiner_m_axis_tvalid; // @[BFS.scala 666:26]
  wire  combiner_m_axis_tready; // @[BFS.scala 666:26]
  wire  combiner_m_axis_tid; // @[BFS.scala 666:26]
  wire [255:0] combiner_io_s_axis_tdata_lo = {io_ddr_in_1_bits_tdata,io_ddr_in_0_bits_tdata}; // @[BFS.scala 669:98]
  wire [255:0] combiner_io_s_axis_tdata_hi = {io_ddr_in_3_bits_tdata,io_ddr_in_2_bits_tdata}; // @[BFS.scala 669:98]
  wire  _combiner_io_s_axis_tkeep_T_4 = io_ddr_in_0_bits_tkeep[0] & io_ddr_in_0_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_5 = io_ddr_in_0_bits_tkeep[1] & io_ddr_in_0_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_6 = io_ddr_in_0_bits_tkeep[2] & io_ddr_in_0_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_7 = io_ddr_in_0_bits_tkeep[3] & io_ddr_in_0_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_12 = io_ddr_in_1_bits_tkeep[0] & io_ddr_in_1_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_13 = io_ddr_in_1_bits_tkeep[1] & io_ddr_in_1_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_14 = io_ddr_in_1_bits_tkeep[2] & io_ddr_in_1_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_15 = io_ddr_in_1_bits_tkeep[3] & io_ddr_in_1_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_20 = io_ddr_in_2_bits_tkeep[0] & io_ddr_in_2_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_21 = io_ddr_in_2_bits_tkeep[1] & io_ddr_in_2_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_22 = io_ddr_in_2_bits_tkeep[2] & io_ddr_in_2_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_23 = io_ddr_in_2_bits_tkeep[3] & io_ddr_in_2_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_28 = io_ddr_in_3_bits_tkeep[0] & io_ddr_in_3_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_29 = io_ddr_in_3_bits_tkeep[1] & io_ddr_in_3_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_30 = io_ddr_in_3_bits_tkeep[2] & io_ddr_in_3_valid; // @[BFS.scala 670:120]
  wire  _combiner_io_s_axis_tkeep_T_31 = io_ddr_in_3_bits_tkeep[3] & io_ddr_in_3_valid; // @[BFS.scala 670:120]
  wire [7:0] combiner_io_s_axis_tkeep_lo = {_combiner_io_s_axis_tkeep_T_15,_combiner_io_s_axis_tkeep_T_14,
    _combiner_io_s_axis_tkeep_T_13,_combiner_io_s_axis_tkeep_T_12,_combiner_io_s_axis_tkeep_T_7,
    _combiner_io_s_axis_tkeep_T_6,_combiner_io_s_axis_tkeep_T_5,_combiner_io_s_axis_tkeep_T_4}; // @[BFS.scala 670:150]
  wire [15:0] _combiner_io_s_axis_tkeep_T_32 = {_combiner_io_s_axis_tkeep_T_31,_combiner_io_s_axis_tkeep_T_30,
    _combiner_io_s_axis_tkeep_T_29,_combiner_io_s_axis_tkeep_T_28,_combiner_io_s_axis_tkeep_T_23,
    _combiner_io_s_axis_tkeep_T_22,_combiner_io_s_axis_tkeep_T_21,_combiner_io_s_axis_tkeep_T_20,
    combiner_io_s_axis_tkeep_lo}; // @[BFS.scala 670:150]
  wire  _combiner_io_s_axis_tvalid_T_2 = io_ddr_in_0_valid | io_ddr_in_1_valid | io_ddr_in_2_valid | io_ddr_in_3_valid; // @[BFS.scala 672:99]
  wire [1:0] combiner_io_s_axis_tvalid_lo = {_combiner_io_s_axis_tvalid_T_2,_combiner_io_s_axis_tvalid_T_2}; // @[BFS.scala 672:111]
  wire [7:0] xbar_io_m_axis_tready_lo = {io_pe_out_7_ready,io_pe_out_6_ready,io_pe_out_5_ready,io_pe_out_4_ready,
    io_pe_out_3_ready,io_pe_out_2_ready,io_pe_out_1_ready,io_pe_out_0_ready}; // @[BFS.scala 689:12]
  wire [7:0] xbar_io_m_axis_tready_hi = {io_pe_out_15_ready,io_pe_out_14_ready,io_pe_out_13_ready,io_pe_out_12_ready,
    io_pe_out_11_ready,io_pe_out_10_ready,io_pe_out_9_ready,io_pe_out_8_ready}; // @[BFS.scala 689:12]
  axis_broadcaster xbar ( // @[BFS.scala 660:20]
    .aclk(xbar_aclk),
    .aresetn(xbar_aresetn),
    .s_axis_tdata(xbar_s_axis_tdata),
    .s_axis_tkeep(xbar_s_axis_tkeep),
    .s_axis_tlast(xbar_s_axis_tlast),
    .s_axis_tvalid(xbar_s_axis_tvalid),
    .s_axis_tready(xbar_s_axis_tready),
    .s_axis_tid(xbar_s_axis_tid),
    .m_axis_tdata(xbar_m_axis_tdata),
    .m_axis_tkeep(xbar_m_axis_tkeep),
    .m_axis_tlast(xbar_m_axis_tlast),
    .m_axis_tvalid(xbar_m_axis_tvalid),
    .m_axis_tready(xbar_m_axis_tready),
    .m_axis_tid(xbar_m_axis_tid)
  );
  axis_combiner combiner ( // @[BFS.scala 666:26]
    .aclk(combiner_aclk),
    .aresetn(combiner_aresetn),
    .s_axis_tdata(combiner_s_axis_tdata),
    .s_axis_tkeep(combiner_s_axis_tkeep),
    .s_axis_tlast(combiner_s_axis_tlast),
    .s_axis_tvalid(combiner_s_axis_tvalid),
    .s_axis_tready(combiner_s_axis_tready),
    .s_axis_tid(combiner_s_axis_tid),
    .m_axis_tdata(combiner_m_axis_tdata),
    .m_axis_tkeep(combiner_m_axis_tkeep),
    .m_axis_tlast(combiner_m_axis_tlast),
    .m_axis_tvalid(combiner_m_axis_tvalid),
    .m_axis_tready(combiner_m_axis_tready),
    .m_axis_tid(combiner_m_axis_tid)
  );
  assign io_ddr_in_0_ready = combiner_s_axis_tready[0]; // @[BFS.scala 674:60]
  assign io_ddr_in_1_ready = combiner_s_axis_tready[1]; // @[BFS.scala 674:60]
  assign io_ddr_in_2_ready = combiner_s_axis_tready[2]; // @[BFS.scala 674:60]
  assign io_ddr_in_3_ready = combiner_s_axis_tready[3]; // @[BFS.scala 674:60]
  assign io_pe_out_0_valid = xbar_m_axis_tvalid[0]; // @[BFS.scala 684:40]
  assign io_pe_out_0_bits_tdata = xbar_m_axis_tdata[511:0]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_0_bits_tkeep = xbar_m_axis_tkeep[15:0]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_1_valid = xbar_m_axis_tvalid[1]; // @[BFS.scala 684:40]
  assign io_pe_out_1_bits_tdata = xbar_m_axis_tdata[1023:512]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_1_bits_tkeep = xbar_m_axis_tkeep[79:64]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_2_valid = xbar_m_axis_tvalid[2]; // @[BFS.scala 684:40]
  assign io_pe_out_2_bits_tdata = xbar_m_axis_tdata[1535:1024]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_2_bits_tkeep = xbar_m_axis_tkeep[143:128]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_3_valid = xbar_m_axis_tvalid[3]; // @[BFS.scala 684:40]
  assign io_pe_out_3_bits_tdata = xbar_m_axis_tdata[2047:1536]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_3_bits_tkeep = xbar_m_axis_tkeep[207:192]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_4_valid = xbar_m_axis_tvalid[4]; // @[BFS.scala 684:40]
  assign io_pe_out_4_bits_tdata = xbar_m_axis_tdata[2559:2048]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_4_bits_tkeep = xbar_m_axis_tkeep[271:256]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_5_valid = xbar_m_axis_tvalid[5]; // @[BFS.scala 684:40]
  assign io_pe_out_5_bits_tdata = xbar_m_axis_tdata[3071:2560]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_5_bits_tkeep = xbar_m_axis_tkeep[335:320]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_6_valid = xbar_m_axis_tvalid[6]; // @[BFS.scala 684:40]
  assign io_pe_out_6_bits_tdata = xbar_m_axis_tdata[3583:3072]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_6_bits_tkeep = xbar_m_axis_tkeep[399:384]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_7_valid = xbar_m_axis_tvalid[7]; // @[BFS.scala 684:40]
  assign io_pe_out_7_bits_tdata = xbar_m_axis_tdata[4095:3584]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_7_bits_tkeep = xbar_m_axis_tkeep[463:448]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_8_valid = xbar_m_axis_tvalid[8]; // @[BFS.scala 684:40]
  assign io_pe_out_8_bits_tdata = xbar_m_axis_tdata[4607:4096]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_8_bits_tkeep = xbar_m_axis_tkeep[527:512]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_9_valid = xbar_m_axis_tvalid[9]; // @[BFS.scala 684:40]
  assign io_pe_out_9_bits_tdata = xbar_m_axis_tdata[5119:4608]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_9_bits_tkeep = xbar_m_axis_tkeep[591:576]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_10_valid = xbar_m_axis_tvalid[10]; // @[BFS.scala 684:40]
  assign io_pe_out_10_bits_tdata = xbar_m_axis_tdata[5631:5120]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_10_bits_tkeep = xbar_m_axis_tkeep[655:640]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_11_valid = xbar_m_axis_tvalid[11]; // @[BFS.scala 684:40]
  assign io_pe_out_11_bits_tdata = xbar_m_axis_tdata[6143:5632]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_11_bits_tkeep = xbar_m_axis_tkeep[719:704]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_12_valid = xbar_m_axis_tvalid[12]; // @[BFS.scala 684:40]
  assign io_pe_out_12_bits_tdata = xbar_m_axis_tdata[6655:6144]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_12_bits_tkeep = xbar_m_axis_tkeep[783:768]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_13_valid = xbar_m_axis_tvalid[13]; // @[BFS.scala 684:40]
  assign io_pe_out_13_bits_tdata = xbar_m_axis_tdata[7167:6656]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_13_bits_tkeep = xbar_m_axis_tkeep[847:832]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_14_valid = xbar_m_axis_tvalid[14]; // @[BFS.scala 684:40]
  assign io_pe_out_14_bits_tdata = xbar_m_axis_tdata[7679:7168]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_14_bits_tkeep = xbar_m_axis_tkeep[911:896]; // @[nf_arm_doce_top.scala 113:13]
  assign io_pe_out_15_valid = xbar_m_axis_tvalid[15]; // @[BFS.scala 684:40]
  assign io_pe_out_15_bits_tdata = xbar_m_axis_tdata[8191:7680]; // @[nf_arm_doce_top.scala 111:21]
  assign io_pe_out_15_bits_tkeep = xbar_m_axis_tkeep[975:960]; // @[nf_arm_doce_top.scala 113:13]
  assign xbar_aclk = clock; // @[BFS.scala 679:31]
  assign xbar_aresetn = ~reset; // @[BFS.scala 680:22]
  assign xbar_s_axis_tdata = combiner_m_axis_tdata; // @[BFS.scala 676:20]
  assign xbar_s_axis_tkeep = combiner_m_axis_tkeep; // @[BFS.scala 676:20]
  assign xbar_s_axis_tlast = combiner_m_axis_tlast; // @[BFS.scala 676:20]
  assign xbar_s_axis_tvalid = combiner_m_axis_tvalid; // @[BFS.scala 676:20]
  assign xbar_s_axis_tid = combiner_m_axis_tid; // @[BFS.scala 676:20]
  assign xbar_m_axis_tready = {xbar_io_m_axis_tready_hi,xbar_io_m_axis_tready_lo}; // @[BFS.scala 689:12]
  assign combiner_aclk = clock; // @[BFS.scala 667:37]
  assign combiner_aresetn = ~reset; // @[BFS.scala 668:28]
  assign combiner_s_axis_tdata = {combiner_io_s_axis_tdata_hi,combiner_io_s_axis_tdata_lo}; // @[BFS.scala 669:98]
  assign combiner_s_axis_tkeep = {{48'd0}, _combiner_io_s_axis_tkeep_T_32}; // @[BFS.scala 670:150]
  assign combiner_s_axis_tlast = 4'hf; // @[BFS.scala 671:98]
  assign combiner_s_axis_tvalid = {combiner_io_s_axis_tvalid_lo,combiner_io_s_axis_tvalid_lo}; // @[BFS.scala 672:111]
  assign combiner_s_axis_tid = 4'h0;
  assign combiner_m_axis_tready = xbar_s_axis_tready; // @[BFS.scala 676:20]
endmodule
module BFS_ps(
  input          clock,
  input          reset,
  input  [63:0]  io_config_awaddr,
  input          io_config_awvalid,
  output         io_config_awready,
  input  [63:0]  io_config_araddr,
  input          io_config_arvalid,
  output         io_config_arready,
  input  [31:0]  io_config_wdata,
  input  [3:0]   io_config_wstrb,
  input          io_config_wvalid,
  output         io_config_wready,
  output [31:0]  io_config_rdata,
  output [1:0]   io_config_rresp,
  output         io_config_rvalid,
  input          io_config_rready,
  output [1:0]   io_config_bresp,
  output         io_config_bvalid,
  input          io_config_bready,
  input          io_PLmemory_0_aw_ready,
  output         io_PLmemory_0_aw_valid,
  output [63:0]  io_PLmemory_0_aw_bits_awaddr,
  output [6:0]   io_PLmemory_0_aw_bits_awid,
  output [7:0]   io_PLmemory_0_aw_bits_awlen,
  output [2:0]   io_PLmemory_0_aw_bits_awsize,
  output [1:0]   io_PLmemory_0_aw_bits_awburst,
  output         io_PLmemory_0_aw_bits_awlock,
  input          io_PLmemory_0_ar_ready,
  output         io_PLmemory_0_ar_valid,
  output [63:0]  io_PLmemory_0_ar_bits_araddr,
  output [6:0]   io_PLmemory_0_ar_bits_arid,
  output [7:0]   io_PLmemory_0_ar_bits_arlen,
  output [2:0]   io_PLmemory_0_ar_bits_arsize,
  output [1:0]   io_PLmemory_0_ar_bits_arburst,
  output         io_PLmemory_0_ar_bits_arlock,
  input          io_PLmemory_0_w_ready,
  output         io_PLmemory_0_w_valid,
  output [511:0] io_PLmemory_0_w_bits_wdata,
  output [63:0]  io_PLmemory_0_w_bits_wstrb,
  output         io_PLmemory_0_w_bits_wlast,
  output         io_PLmemory_0_r_ready,
  input          io_PLmemory_0_r_valid,
  input  [511:0] io_PLmemory_0_r_bits_rdata,
  input  [6:0]   io_PLmemory_0_r_bits_rid,
  input          io_PLmemory_0_r_bits_rlast,
  output         io_PLmemory_0_b_ready,
  input          io_PLmemory_0_b_valid,
  input  [1:0]   io_PLmemory_0_b_bits_bresp,
  input  [6:0]   io_PLmemory_0_b_bits_bid,
  input          io_PLmemory_1_aw_ready,
  output         io_PLmemory_1_aw_valid,
  output [63:0]  io_PLmemory_1_aw_bits_awaddr,
  output [6:0]   io_PLmemory_1_aw_bits_awid,
  output [7:0]   io_PLmemory_1_aw_bits_awlen,
  output [2:0]   io_PLmemory_1_aw_bits_awsize,
  output [1:0]   io_PLmemory_1_aw_bits_awburst,
  output         io_PLmemory_1_aw_bits_awlock,
  input          io_PLmemory_1_ar_ready,
  output         io_PLmemory_1_ar_valid,
  output [63:0]  io_PLmemory_1_ar_bits_araddr,
  output [6:0]   io_PLmemory_1_ar_bits_arid,
  output [7:0]   io_PLmemory_1_ar_bits_arlen,
  output [2:0]   io_PLmemory_1_ar_bits_arsize,
  output [1:0]   io_PLmemory_1_ar_bits_arburst,
  output         io_PLmemory_1_ar_bits_arlock,
  input          io_PLmemory_1_w_ready,
  output         io_PLmemory_1_w_valid,
  output [511:0] io_PLmemory_1_w_bits_wdata,
  output [63:0]  io_PLmemory_1_w_bits_wstrb,
  output         io_PLmemory_1_w_bits_wlast,
  output         io_PLmemory_1_r_ready,
  input          io_PLmemory_1_r_valid,
  input  [511:0] io_PLmemory_1_r_bits_rdata,
  input  [6:0]   io_PLmemory_1_r_bits_rid,
  input          io_PLmemory_1_r_bits_rlast,
  output         io_PLmemory_1_b_ready,
  input          io_PLmemory_1_b_valid,
  input  [1:0]   io_PLmemory_1_b_bits_bresp,
  input  [6:0]   io_PLmemory_1_b_bits_bid,
  input          io_PSmemory_0_aw_ready,
  output         io_PSmemory_0_aw_valid,
  output [63:0]  io_PSmemory_0_aw_bits_awaddr,
  output [5:0]   io_PSmemory_0_aw_bits_awid,
  output [7:0]   io_PSmemory_0_aw_bits_awlen,
  output [2:0]   io_PSmemory_0_aw_bits_awsize,
  output [1:0]   io_PSmemory_0_aw_bits_awburst,
  output         io_PSmemory_0_aw_bits_awlock,
  input          io_PSmemory_0_ar_ready,
  output         io_PSmemory_0_ar_valid,
  output [63:0]  io_PSmemory_0_ar_bits_araddr,
  output [5:0]   io_PSmemory_0_ar_bits_arid,
  output [7:0]   io_PSmemory_0_ar_bits_arlen,
  output [2:0]   io_PSmemory_0_ar_bits_arsize,
  output [1:0]   io_PSmemory_0_ar_bits_arburst,
  output         io_PSmemory_0_ar_bits_arlock,
  input          io_PSmemory_0_w_ready,
  output         io_PSmemory_0_w_valid,
  output [127:0] io_PSmemory_0_w_bits_wdata,
  output [15:0]  io_PSmemory_0_w_bits_wstrb,
  output         io_PSmemory_0_w_bits_wlast,
  output         io_PSmemory_0_r_ready,
  input          io_PSmemory_0_r_valid,
  input  [127:0] io_PSmemory_0_r_bits_rdata,
  input  [5:0]   io_PSmemory_0_r_bits_rid,
  input          io_PSmemory_0_r_bits_rlast,
  output         io_PSmemory_0_b_ready,
  input          io_PSmemory_0_b_valid,
  input  [1:0]   io_PSmemory_0_b_bits_bresp,
  input  [5:0]   io_PSmemory_0_b_bits_bid,
  input          io_PSmemory_1_aw_ready,
  output         io_PSmemory_1_aw_valid,
  output [63:0]  io_PSmemory_1_aw_bits_awaddr,
  output [5:0]   io_PSmemory_1_aw_bits_awid,
  output [7:0]   io_PSmemory_1_aw_bits_awlen,
  output [2:0]   io_PSmemory_1_aw_bits_awsize,
  output [1:0]   io_PSmemory_1_aw_bits_awburst,
  output         io_PSmemory_1_aw_bits_awlock,
  input          io_PSmemory_1_ar_ready,
  output         io_PSmemory_1_ar_valid,
  output [63:0]  io_PSmemory_1_ar_bits_araddr,
  output [5:0]   io_PSmemory_1_ar_bits_arid,
  output [7:0]   io_PSmemory_1_ar_bits_arlen,
  output [2:0]   io_PSmemory_1_ar_bits_arsize,
  output [1:0]   io_PSmemory_1_ar_bits_arburst,
  output         io_PSmemory_1_ar_bits_arlock,
  input          io_PSmemory_1_w_ready,
  output         io_PSmemory_1_w_valid,
  output [127:0] io_PSmemory_1_w_bits_wdata,
  output [15:0]  io_PSmemory_1_w_bits_wstrb,
  output         io_PSmemory_1_w_bits_wlast,
  output         io_PSmemory_1_r_ready,
  input          io_PSmemory_1_r_valid,
  input  [127:0] io_PSmemory_1_r_bits_rdata,
  input  [5:0]   io_PSmemory_1_r_bits_rid,
  input          io_PSmemory_1_r_bits_rlast,
  output         io_PSmemory_1_b_ready,
  input          io_PSmemory_1_b_valid,
  input  [1:0]   io_PSmemory_1_b_bits_bresp,
  input  [5:0]   io_PSmemory_1_b_bits_bid,
  input          io_PSmemory_2_aw_ready,
  output         io_PSmemory_2_aw_valid,
  output [63:0]  io_PSmemory_2_aw_bits_awaddr,
  output [5:0]   io_PSmemory_2_aw_bits_awid,
  output [7:0]   io_PSmemory_2_aw_bits_awlen,
  output [2:0]   io_PSmemory_2_aw_bits_awsize,
  output [1:0]   io_PSmemory_2_aw_bits_awburst,
  output         io_PSmemory_2_aw_bits_awlock,
  input          io_PSmemory_2_ar_ready,
  output         io_PSmemory_2_ar_valid,
  output [63:0]  io_PSmemory_2_ar_bits_araddr,
  output [5:0]   io_PSmemory_2_ar_bits_arid,
  output [7:0]   io_PSmemory_2_ar_bits_arlen,
  output [2:0]   io_PSmemory_2_ar_bits_arsize,
  output [1:0]   io_PSmemory_2_ar_bits_arburst,
  output         io_PSmemory_2_ar_bits_arlock,
  input          io_PSmemory_2_w_ready,
  output         io_PSmemory_2_w_valid,
  output [127:0] io_PSmemory_2_w_bits_wdata,
  output [15:0]  io_PSmemory_2_w_bits_wstrb,
  output         io_PSmemory_2_w_bits_wlast,
  output         io_PSmemory_2_r_ready,
  input          io_PSmemory_2_r_valid,
  input  [127:0] io_PSmemory_2_r_bits_rdata,
  input  [5:0]   io_PSmemory_2_r_bits_rid,
  input          io_PSmemory_2_r_bits_rlast,
  output         io_PSmemory_2_b_ready,
  input          io_PSmemory_2_b_valid,
  input  [1:0]   io_PSmemory_2_b_bits_bresp,
  input  [5:0]   io_PSmemory_2_b_bits_bid,
  input          io_PSmemory_3_aw_ready,
  output         io_PSmemory_3_aw_valid,
  output [63:0]  io_PSmemory_3_aw_bits_awaddr,
  output [5:0]   io_PSmemory_3_aw_bits_awid,
  output [7:0]   io_PSmemory_3_aw_bits_awlen,
  output [2:0]   io_PSmemory_3_aw_bits_awsize,
  output [1:0]   io_PSmemory_3_aw_bits_awburst,
  output         io_PSmemory_3_aw_bits_awlock,
  input          io_PSmemory_3_ar_ready,
  output         io_PSmemory_3_ar_valid,
  output [63:0]  io_PSmemory_3_ar_bits_araddr,
  output [5:0]   io_PSmemory_3_ar_bits_arid,
  output [7:0]   io_PSmemory_3_ar_bits_arlen,
  output [2:0]   io_PSmemory_3_ar_bits_arsize,
  output [1:0]   io_PSmemory_3_ar_bits_arburst,
  output         io_PSmemory_3_ar_bits_arlock,
  input          io_PSmemory_3_w_ready,
  output         io_PSmemory_3_w_valid,
  output [127:0] io_PSmemory_3_w_bits_wdata,
  output [15:0]  io_PSmemory_3_w_bits_wstrb,
  output         io_PSmemory_3_w_bits_wlast,
  output         io_PSmemory_3_r_ready,
  input          io_PSmemory_3_r_valid,
  input  [127:0] io_PSmemory_3_r_bits_rdata,
  input  [5:0]   io_PSmemory_3_r_bits_rid,
  input          io_PSmemory_3_r_bits_rlast,
  output         io_PSmemory_3_b_ready,
  input          io_PSmemory_3_b_valid,
  input  [1:0]   io_PSmemory_3_b_bits_bresp,
  input  [5:0]   io_PSmemory_3_b_bits_bid
);
  wire  controls_clock; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_reset; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_0; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_1; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_2; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_3; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_4; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_5; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_6; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_7; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_8; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_9; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_10; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_data_11; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_0; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_1; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_2; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_3; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_4; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_5; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_6; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_7; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_8; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_9; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_10; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_11; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_12; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_13; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_14; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_fin_15; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_signal; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_start; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_level; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_unvisited_size; // @[nf_arm_doce_top_main.scala 31:24]
  wire [63:0] controls_io_traveled_edges; // @[nf_arm_doce_top_main.scala 31:24]
  wire [63:0] controls_io_config_awaddr; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_config_awready; // @[nf_arm_doce_top_main.scala 31:24]
  wire [63:0] controls_io_config_araddr; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_config_arvalid; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_config_arready; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_config_wdata; // @[nf_arm_doce_top_main.scala 31:24]
  wire [3:0] controls_io_config_wstrb; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_config_wvalid; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_config_wready; // @[nf_arm_doce_top_main.scala 31:24]
  wire [31:0] controls_io_config_rdata; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_config_rvalid; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_config_rready; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_config_bvalid; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_config_bready; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_flush_cache; // @[nf_arm_doce_top_main.scala 31:24]
  wire  controls_io_flush_cache_end; // @[nf_arm_doce_top_main.scala 31:24]
  wire  pl_mc_clock; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_reset; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_out_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_out_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [511:0] pl_mc_io_cacheable_out_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire [15:0] pl_mc_io_cacheable_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_0_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_0_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_0_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_1_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_1_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_1_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_2_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_2_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_2_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_3_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_3_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_3_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_4_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_4_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_4_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_5_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_5_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_5_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_6_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_6_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_6_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_7_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_7_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_7_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_8_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_8_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_8_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_9_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_9_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_9_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_10_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_10_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_10_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_11_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_11_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_11_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_12_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_12_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_12_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_13_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_13_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_13_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_14_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_14_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_14_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_15_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_cacheable_in_15_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_cacheable_in_15_bits_tdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_non_cacheable_in_aw_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_non_cacheable_in_aw_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [63:0] pl_mc_io_non_cacheable_in_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 33:21]
  wire [6:0] pl_mc_io_non_cacheable_in_aw_bits_awid; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_non_cacheable_in_w_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_non_cacheable_in_w_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [511:0] pl_mc_io_non_cacheable_in_w_bits_wdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire [63:0] pl_mc_io_non_cacheable_in_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_0_aw_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_0_aw_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [63:0] pl_mc_io_ddr_out_0_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_0_ar_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_0_ar_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [63:0] pl_mc_io_ddr_out_0_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_0_w_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_0_w_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [511:0] pl_mc_io_ddr_out_0_w_bits_wdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_0_w_bits_wlast; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_0_r_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [511:0] pl_mc_io_ddr_out_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_1_aw_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_1_aw_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [63:0] pl_mc_io_ddr_out_1_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 33:21]
  wire [6:0] pl_mc_io_ddr_out_1_aw_bits_awid; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_1_w_ready; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_ddr_out_1_w_valid; // @[nf_arm_doce_top_main.scala 33:21]
  wire [511:0] pl_mc_io_ddr_out_1_w_bits_wdata; // @[nf_arm_doce_top_main.scala 33:21]
  wire [63:0] pl_mc_io_ddr_out_1_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 33:21]
  wire [63:0] pl_mc_io_tiers_base_addr_0; // @[nf_arm_doce_top_main.scala 33:21]
  wire [63:0] pl_mc_io_tiers_base_addr_1; // @[nf_arm_doce_top_main.scala 33:21]
  wire [31:0] pl_mc_io_unvisited_size; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_start; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_signal; // @[nf_arm_doce_top_main.scala 33:21]
  wire  pl_mc_io_end; // @[nf_arm_doce_top_main.scala 33:21]
  wire  Scatters_0_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_0_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_0_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_0_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_0_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_0_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_0_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_0_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_0_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_1_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_1_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_1_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_1_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_1_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_1_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_1_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_1_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_1_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_2_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_2_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_2_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_2_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_2_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_2_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_2_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_2_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_2_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_3_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_3_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_3_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_3_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_3_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_3_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_3_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_3_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_3_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_4_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_4_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_4_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_4_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_4_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_4_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_4_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_4_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_4_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_4_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_5_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_5_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_5_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_5_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_5_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_5_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_5_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_5_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_5_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_5_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_6_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_6_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_6_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_6_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_6_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_6_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_6_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_6_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_6_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_6_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_7_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_7_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_7_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_7_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_7_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_7_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_7_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_7_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_7_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_7_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_8_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_8_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_8_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_8_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_8_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_8_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_8_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_8_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_8_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_8_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_9_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_9_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_9_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_9_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_9_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_9_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_9_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_9_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_9_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_9_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_10_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_10_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_10_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_10_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_10_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_10_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_10_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_10_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_10_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_10_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_11_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_11_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_11_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_11_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_11_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_11_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_11_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_11_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_11_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_11_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_12_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_12_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_12_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_12_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_12_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_12_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_12_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_12_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_12_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_12_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_13_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_13_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_13_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_13_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_13_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_13_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_13_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_13_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_13_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_13_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_14_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_14_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_14_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_14_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_14_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_14_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_14_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_14_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_14_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_14_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_15_clock; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_15_reset; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_15_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_15_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [511:0] Scatters_15_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire [15:0] Scatters_15_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_15_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_15_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 35:16]
  wire [31:0] Scatters_15_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Scatters_15_io_end; // @[nf_arm_doce_top_main.scala 35:16]
  wire  Gathers_clock; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_reset; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_ddr_in_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_ddr_in_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [511:0] Gathers_io_ddr_in_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire [15:0] Gathers_io_ddr_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_0_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_0_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [31:0] Gathers_io_gather_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_1_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_1_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [31:0] Gathers_io_gather_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_2_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_2_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [31:0] Gathers_io_gather_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_3_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_3_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [31:0] Gathers_io_gather_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_4_ready; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Gathers_io_gather_out_4_valid; // @[nf_arm_doce_top_main.scala 37:23]
  wire [31:0] Gathers_io_gather_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 37:23]
  wire  Applys_clock; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Applys_reset; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Applys_io_ddr_aw_ready; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Applys_io_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 38:22]
  wire [63:0] Applys_io_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 38:22]
  wire [6:0] Applys_io_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Applys_io_ddr_w_ready; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Applys_io_ddr_w_valid; // @[nf_arm_doce_top_main.scala 38:22]
  wire [511:0] Applys_io_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 38:22]
  wire [63:0] Applys_io_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Applys_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Applys_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 38:22]
  wire [31:0] Applys_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 38:22]
  wire [31:0] Applys_io_level; // @[nf_arm_doce_top_main.scala 38:22]
  wire [63:0] Applys_io_level_base_addr; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Applys_io_end; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Applys_io_flush; // @[nf_arm_doce_top_main.scala 38:22]
  wire  Broadcasts_0_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_0_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Broadcasts_0_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [7:0] Broadcasts_0_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 40:16]
  wire [2:0] Broadcasts_0_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Broadcasts_0_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Broadcasts_0_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Broadcasts_0_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Broadcasts_0_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Broadcasts_0_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_0_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_0_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_signal; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_0_io_traveled_edges; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_start; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Broadcasts_0_io_root; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_0_io_issue_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Broadcasts_0_io_recv_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_1_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Broadcasts_1_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [7:0] Broadcasts_1_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 40:16]
  wire [2:0] Broadcasts_1_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Broadcasts_1_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Broadcasts_1_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Broadcasts_1_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Broadcasts_1_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Broadcasts_1_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_1_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_1_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_signal; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_1_io_traveled_edges; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_1_io_issue_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Broadcasts_1_io_recv_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_2_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Broadcasts_2_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [7:0] Broadcasts_2_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 40:16]
  wire [2:0] Broadcasts_2_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Broadcasts_2_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Broadcasts_2_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Broadcasts_2_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Broadcasts_2_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Broadcasts_2_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_2_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_2_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_signal; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_2_io_traveled_edges; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_2_io_issue_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Broadcasts_2_io_recv_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_3_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Broadcasts_3_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [7:0] Broadcasts_3_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 40:16]
  wire [2:0] Broadcasts_3_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Broadcasts_3_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [5:0] Broadcasts_3_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Broadcasts_3_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [127:0] Broadcasts_3_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Broadcasts_3_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_3_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_3_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_signal; // @[nf_arm_doce_top_main.scala 40:16]
  wire [63:0] Broadcasts_3_io_traveled_edges; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Broadcasts_3_io_issue_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire [3:0] Broadcasts_3_io_recv_sync; // @[nf_arm_doce_top_main.scala 40:16]
  wire  bxbar_clock; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_reset; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_ddr_in_0_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_ddr_in_0_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [127:0] bxbar_io_ddr_in_0_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [3:0] bxbar_io_ddr_in_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_ddr_in_1_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_ddr_in_1_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [127:0] bxbar_io_ddr_in_1_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [3:0] bxbar_io_ddr_in_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_ddr_in_2_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_ddr_in_2_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [127:0] bxbar_io_ddr_in_2_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [3:0] bxbar_io_ddr_in_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_ddr_in_3_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_ddr_in_3_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [127:0] bxbar_io_ddr_in_3_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [3:0] bxbar_io_ddr_in_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_0_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_0_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_1_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_1_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_2_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_2_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_3_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_3_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_4_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_4_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_4_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_5_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_5_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_5_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_5_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_6_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_6_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_6_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_6_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_7_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_7_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_7_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_7_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_8_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_8_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_8_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_8_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_9_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_9_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_9_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_9_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_10_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_10_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_10_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_10_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_11_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_11_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_11_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_11_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_12_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_12_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_12_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_12_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_13_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_13_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_13_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_13_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_14_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_14_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_14_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_14_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_15_ready; // @[nf_arm_doce_top_main.scala 43:21]
  wire  bxbar_io_pe_out_15_valid; // @[nf_arm_doce_top_main.scala 43:21]
  wire [511:0] bxbar_io_pe_out_15_bits_tdata; // @[nf_arm_doce_top_main.scala 43:21]
  wire [15:0] bxbar_io_pe_out_15_bits_tkeep; // @[nf_arm_doce_top_main.scala 43:21]
  wire  _Broadcasts_0_io_recv_sync_WIRE_1 = Broadcasts_1_io_issue_sync; // @[nf_arm_doce_top_main.scala 59:32 nf_arm_doce_top_main.scala 59:32]
  wire  _Broadcasts_0_io_recv_sync_WIRE_0 = Broadcasts_0_io_issue_sync; // @[nf_arm_doce_top_main.scala 59:32 nf_arm_doce_top_main.scala 59:32]
  wire [1:0] Broadcasts_0_io_recv_sync_lo = {_Broadcasts_0_io_recv_sync_WIRE_1,_Broadcasts_0_io_recv_sync_WIRE_0}; // @[nf_arm_doce_top_main.scala 59:77]
  wire  _Broadcasts_0_io_recv_sync_WIRE_3 = Broadcasts_3_io_issue_sync; // @[nf_arm_doce_top_main.scala 59:32 nf_arm_doce_top_main.scala 59:32]
  wire  _Broadcasts_0_io_recv_sync_WIRE_2 = Broadcasts_2_io_issue_sync; // @[nf_arm_doce_top_main.scala 59:32 nf_arm_doce_top_main.scala 59:32]
  wire [1:0] Broadcasts_0_io_recv_sync_hi = {_Broadcasts_0_io_recv_sync_WIRE_3,_Broadcasts_0_io_recv_sync_WIRE_2}; // @[nf_arm_doce_top_main.scala 59:77]
  wire [63:0] _controls_io_traveled_edges_T_1 = Broadcasts_0_io_traveled_edges + Broadcasts_1_io_traveled_edges; // @[nf_arm_doce_top_main.scala 91:82]
  wire [63:0] _controls_io_traveled_edges_T_3 = _controls_io_traveled_edges_T_1 + Broadcasts_2_io_traveled_edges; // @[nf_arm_doce_top_main.scala 91:82]
  controller controls ( // @[nf_arm_doce_top_main.scala 31:24]
    .clock(controls_clock),
    .reset(controls_reset),
    .io_data_0(controls_io_data_0),
    .io_data_1(controls_io_data_1),
    .io_data_2(controls_io_data_2),
    .io_data_3(controls_io_data_3),
    .io_data_4(controls_io_data_4),
    .io_data_5(controls_io_data_5),
    .io_data_6(controls_io_data_6),
    .io_data_7(controls_io_data_7),
    .io_data_8(controls_io_data_8),
    .io_data_9(controls_io_data_9),
    .io_data_10(controls_io_data_10),
    .io_data_11(controls_io_data_11),
    .io_fin_0(controls_io_fin_0),
    .io_fin_1(controls_io_fin_1),
    .io_fin_2(controls_io_fin_2),
    .io_fin_3(controls_io_fin_3),
    .io_fin_4(controls_io_fin_4),
    .io_fin_5(controls_io_fin_5),
    .io_fin_6(controls_io_fin_6),
    .io_fin_7(controls_io_fin_7),
    .io_fin_8(controls_io_fin_8),
    .io_fin_9(controls_io_fin_9),
    .io_fin_10(controls_io_fin_10),
    .io_fin_11(controls_io_fin_11),
    .io_fin_12(controls_io_fin_12),
    .io_fin_13(controls_io_fin_13),
    .io_fin_14(controls_io_fin_14),
    .io_fin_15(controls_io_fin_15),
    .io_signal(controls_io_signal),
    .io_start(controls_io_start),
    .io_level(controls_io_level),
    .io_unvisited_size(controls_io_unvisited_size),
    .io_traveled_edges(controls_io_traveled_edges),
    .io_config_awaddr(controls_io_config_awaddr),
    .io_config_awready(controls_io_config_awready),
    .io_config_araddr(controls_io_config_araddr),
    .io_config_arvalid(controls_io_config_arvalid),
    .io_config_arready(controls_io_config_arready),
    .io_config_wdata(controls_io_config_wdata),
    .io_config_wstrb(controls_io_config_wstrb),
    .io_config_wvalid(controls_io_config_wvalid),
    .io_config_wready(controls_io_config_wready),
    .io_config_rdata(controls_io_config_rdata),
    .io_config_rvalid(controls_io_config_rvalid),
    .io_config_rready(controls_io_config_rready),
    .io_config_bvalid(controls_io_config_bvalid),
    .io_config_bready(controls_io_config_bready),
    .io_flush_cache(controls_io_flush_cache),
    .io_flush_cache_end(controls_io_flush_cache_end)
  );
  multi_port_mc pl_mc ( // @[nf_arm_doce_top_main.scala 33:21]
    .clock(pl_mc_clock),
    .reset(pl_mc_reset),
    .io_cacheable_out_ready(pl_mc_io_cacheable_out_ready),
    .io_cacheable_out_valid(pl_mc_io_cacheable_out_valid),
    .io_cacheable_out_bits_tdata(pl_mc_io_cacheable_out_bits_tdata),
    .io_cacheable_out_bits_tkeep(pl_mc_io_cacheable_out_bits_tkeep),
    .io_cacheable_in_0_ready(pl_mc_io_cacheable_in_0_ready),
    .io_cacheable_in_0_valid(pl_mc_io_cacheable_in_0_valid),
    .io_cacheable_in_0_bits_tdata(pl_mc_io_cacheable_in_0_bits_tdata),
    .io_cacheable_in_1_ready(pl_mc_io_cacheable_in_1_ready),
    .io_cacheable_in_1_valid(pl_mc_io_cacheable_in_1_valid),
    .io_cacheable_in_1_bits_tdata(pl_mc_io_cacheable_in_1_bits_tdata),
    .io_cacheable_in_2_ready(pl_mc_io_cacheable_in_2_ready),
    .io_cacheable_in_2_valid(pl_mc_io_cacheable_in_2_valid),
    .io_cacheable_in_2_bits_tdata(pl_mc_io_cacheable_in_2_bits_tdata),
    .io_cacheable_in_3_ready(pl_mc_io_cacheable_in_3_ready),
    .io_cacheable_in_3_valid(pl_mc_io_cacheable_in_3_valid),
    .io_cacheable_in_3_bits_tdata(pl_mc_io_cacheable_in_3_bits_tdata),
    .io_cacheable_in_4_ready(pl_mc_io_cacheable_in_4_ready),
    .io_cacheable_in_4_valid(pl_mc_io_cacheable_in_4_valid),
    .io_cacheable_in_4_bits_tdata(pl_mc_io_cacheable_in_4_bits_tdata),
    .io_cacheable_in_5_ready(pl_mc_io_cacheable_in_5_ready),
    .io_cacheable_in_5_valid(pl_mc_io_cacheable_in_5_valid),
    .io_cacheable_in_5_bits_tdata(pl_mc_io_cacheable_in_5_bits_tdata),
    .io_cacheable_in_6_ready(pl_mc_io_cacheable_in_6_ready),
    .io_cacheable_in_6_valid(pl_mc_io_cacheable_in_6_valid),
    .io_cacheable_in_6_bits_tdata(pl_mc_io_cacheable_in_6_bits_tdata),
    .io_cacheable_in_7_ready(pl_mc_io_cacheable_in_7_ready),
    .io_cacheable_in_7_valid(pl_mc_io_cacheable_in_7_valid),
    .io_cacheable_in_7_bits_tdata(pl_mc_io_cacheable_in_7_bits_tdata),
    .io_cacheable_in_8_ready(pl_mc_io_cacheable_in_8_ready),
    .io_cacheable_in_8_valid(pl_mc_io_cacheable_in_8_valid),
    .io_cacheable_in_8_bits_tdata(pl_mc_io_cacheable_in_8_bits_tdata),
    .io_cacheable_in_9_ready(pl_mc_io_cacheable_in_9_ready),
    .io_cacheable_in_9_valid(pl_mc_io_cacheable_in_9_valid),
    .io_cacheable_in_9_bits_tdata(pl_mc_io_cacheable_in_9_bits_tdata),
    .io_cacheable_in_10_ready(pl_mc_io_cacheable_in_10_ready),
    .io_cacheable_in_10_valid(pl_mc_io_cacheable_in_10_valid),
    .io_cacheable_in_10_bits_tdata(pl_mc_io_cacheable_in_10_bits_tdata),
    .io_cacheable_in_11_ready(pl_mc_io_cacheable_in_11_ready),
    .io_cacheable_in_11_valid(pl_mc_io_cacheable_in_11_valid),
    .io_cacheable_in_11_bits_tdata(pl_mc_io_cacheable_in_11_bits_tdata),
    .io_cacheable_in_12_ready(pl_mc_io_cacheable_in_12_ready),
    .io_cacheable_in_12_valid(pl_mc_io_cacheable_in_12_valid),
    .io_cacheable_in_12_bits_tdata(pl_mc_io_cacheable_in_12_bits_tdata),
    .io_cacheable_in_13_ready(pl_mc_io_cacheable_in_13_ready),
    .io_cacheable_in_13_valid(pl_mc_io_cacheable_in_13_valid),
    .io_cacheable_in_13_bits_tdata(pl_mc_io_cacheable_in_13_bits_tdata),
    .io_cacheable_in_14_ready(pl_mc_io_cacheable_in_14_ready),
    .io_cacheable_in_14_valid(pl_mc_io_cacheable_in_14_valid),
    .io_cacheable_in_14_bits_tdata(pl_mc_io_cacheable_in_14_bits_tdata),
    .io_cacheable_in_15_ready(pl_mc_io_cacheable_in_15_ready),
    .io_cacheable_in_15_valid(pl_mc_io_cacheable_in_15_valid),
    .io_cacheable_in_15_bits_tdata(pl_mc_io_cacheable_in_15_bits_tdata),
    .io_non_cacheable_in_aw_ready(pl_mc_io_non_cacheable_in_aw_ready),
    .io_non_cacheable_in_aw_valid(pl_mc_io_non_cacheable_in_aw_valid),
    .io_non_cacheable_in_aw_bits_awaddr(pl_mc_io_non_cacheable_in_aw_bits_awaddr),
    .io_non_cacheable_in_aw_bits_awid(pl_mc_io_non_cacheable_in_aw_bits_awid),
    .io_non_cacheable_in_w_ready(pl_mc_io_non_cacheable_in_w_ready),
    .io_non_cacheable_in_w_valid(pl_mc_io_non_cacheable_in_w_valid),
    .io_non_cacheable_in_w_bits_wdata(pl_mc_io_non_cacheable_in_w_bits_wdata),
    .io_non_cacheable_in_w_bits_wstrb(pl_mc_io_non_cacheable_in_w_bits_wstrb),
    .io_ddr_out_0_aw_ready(pl_mc_io_ddr_out_0_aw_ready),
    .io_ddr_out_0_aw_valid(pl_mc_io_ddr_out_0_aw_valid),
    .io_ddr_out_0_aw_bits_awaddr(pl_mc_io_ddr_out_0_aw_bits_awaddr),
    .io_ddr_out_0_ar_ready(pl_mc_io_ddr_out_0_ar_ready),
    .io_ddr_out_0_ar_valid(pl_mc_io_ddr_out_0_ar_valid),
    .io_ddr_out_0_ar_bits_araddr(pl_mc_io_ddr_out_0_ar_bits_araddr),
    .io_ddr_out_0_w_ready(pl_mc_io_ddr_out_0_w_ready),
    .io_ddr_out_0_w_valid(pl_mc_io_ddr_out_0_w_valid),
    .io_ddr_out_0_w_bits_wdata(pl_mc_io_ddr_out_0_w_bits_wdata),
    .io_ddr_out_0_w_bits_wlast(pl_mc_io_ddr_out_0_w_bits_wlast),
    .io_ddr_out_0_r_valid(pl_mc_io_ddr_out_0_r_valid),
    .io_ddr_out_0_r_bits_rdata(pl_mc_io_ddr_out_0_r_bits_rdata),
    .io_ddr_out_0_r_bits_rlast(pl_mc_io_ddr_out_0_r_bits_rlast),
    .io_ddr_out_1_aw_ready(pl_mc_io_ddr_out_1_aw_ready),
    .io_ddr_out_1_aw_valid(pl_mc_io_ddr_out_1_aw_valid),
    .io_ddr_out_1_aw_bits_awaddr(pl_mc_io_ddr_out_1_aw_bits_awaddr),
    .io_ddr_out_1_aw_bits_awid(pl_mc_io_ddr_out_1_aw_bits_awid),
    .io_ddr_out_1_w_ready(pl_mc_io_ddr_out_1_w_ready),
    .io_ddr_out_1_w_valid(pl_mc_io_ddr_out_1_w_valid),
    .io_ddr_out_1_w_bits_wdata(pl_mc_io_ddr_out_1_w_bits_wdata),
    .io_ddr_out_1_w_bits_wstrb(pl_mc_io_ddr_out_1_w_bits_wstrb),
    .io_tiers_base_addr_0(pl_mc_io_tiers_base_addr_0),
    .io_tiers_base_addr_1(pl_mc_io_tiers_base_addr_1),
    .io_unvisited_size(pl_mc_io_unvisited_size),
    .io_start(pl_mc_io_start),
    .io_signal(pl_mc_io_signal),
    .io_end(pl_mc_io_end)
  );
  Scatter Scatters_0 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_0_clock),
    .reset(Scatters_0_reset),
    .io_xbar_in_ready(Scatters_0_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_0_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_0_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_0_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_0_io_ddr_out_bits_tdata),
    .io_end(Scatters_0_io_end)
  );
  Scatter_1 Scatters_1 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_1_clock),
    .reset(Scatters_1_reset),
    .io_xbar_in_ready(Scatters_1_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_1_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_1_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_1_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_1_io_ddr_out_bits_tdata),
    .io_end(Scatters_1_io_end)
  );
  Scatter_2 Scatters_2 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_2_clock),
    .reset(Scatters_2_reset),
    .io_xbar_in_ready(Scatters_2_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_2_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_2_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_2_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_2_io_ddr_out_bits_tdata),
    .io_end(Scatters_2_io_end)
  );
  Scatter_3 Scatters_3 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_3_clock),
    .reset(Scatters_3_reset),
    .io_xbar_in_ready(Scatters_3_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_3_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_3_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_3_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_3_io_ddr_out_bits_tdata),
    .io_end(Scatters_3_io_end)
  );
  Scatter_4 Scatters_4 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_4_clock),
    .reset(Scatters_4_reset),
    .io_xbar_in_ready(Scatters_4_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_4_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_4_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_4_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_4_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_4_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_4_io_ddr_out_bits_tdata),
    .io_end(Scatters_4_io_end)
  );
  Scatter_5 Scatters_5 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_5_clock),
    .reset(Scatters_5_reset),
    .io_xbar_in_ready(Scatters_5_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_5_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_5_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_5_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_5_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_5_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_5_io_ddr_out_bits_tdata),
    .io_end(Scatters_5_io_end)
  );
  Scatter_6 Scatters_6 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_6_clock),
    .reset(Scatters_6_reset),
    .io_xbar_in_ready(Scatters_6_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_6_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_6_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_6_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_6_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_6_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_6_io_ddr_out_bits_tdata),
    .io_end(Scatters_6_io_end)
  );
  Scatter_7 Scatters_7 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_7_clock),
    .reset(Scatters_7_reset),
    .io_xbar_in_ready(Scatters_7_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_7_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_7_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_7_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_7_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_7_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_7_io_ddr_out_bits_tdata),
    .io_end(Scatters_7_io_end)
  );
  Scatter_8 Scatters_8 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_8_clock),
    .reset(Scatters_8_reset),
    .io_xbar_in_ready(Scatters_8_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_8_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_8_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_8_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_8_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_8_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_8_io_ddr_out_bits_tdata),
    .io_end(Scatters_8_io_end)
  );
  Scatter_9 Scatters_9 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_9_clock),
    .reset(Scatters_9_reset),
    .io_xbar_in_ready(Scatters_9_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_9_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_9_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_9_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_9_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_9_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_9_io_ddr_out_bits_tdata),
    .io_end(Scatters_9_io_end)
  );
  Scatter_10 Scatters_10 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_10_clock),
    .reset(Scatters_10_reset),
    .io_xbar_in_ready(Scatters_10_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_10_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_10_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_10_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_10_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_10_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_10_io_ddr_out_bits_tdata),
    .io_end(Scatters_10_io_end)
  );
  Scatter_11 Scatters_11 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_11_clock),
    .reset(Scatters_11_reset),
    .io_xbar_in_ready(Scatters_11_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_11_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_11_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_11_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_11_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_11_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_11_io_ddr_out_bits_tdata),
    .io_end(Scatters_11_io_end)
  );
  Scatter_12 Scatters_12 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_12_clock),
    .reset(Scatters_12_reset),
    .io_xbar_in_ready(Scatters_12_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_12_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_12_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_12_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_12_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_12_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_12_io_ddr_out_bits_tdata),
    .io_end(Scatters_12_io_end)
  );
  Scatter_13 Scatters_13 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_13_clock),
    .reset(Scatters_13_reset),
    .io_xbar_in_ready(Scatters_13_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_13_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_13_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_13_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_13_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_13_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_13_io_ddr_out_bits_tdata),
    .io_end(Scatters_13_io_end)
  );
  Scatter_14 Scatters_14 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_14_clock),
    .reset(Scatters_14_reset),
    .io_xbar_in_ready(Scatters_14_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_14_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_14_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_14_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_14_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_14_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_14_io_ddr_out_bits_tdata),
    .io_end(Scatters_14_io_end)
  );
  Scatter_15 Scatters_15 ( // @[nf_arm_doce_top_main.scala 35:16]
    .clock(Scatters_15_clock),
    .reset(Scatters_15_reset),
    .io_xbar_in_ready(Scatters_15_io_xbar_in_ready),
    .io_xbar_in_valid(Scatters_15_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Scatters_15_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Scatters_15_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Scatters_15_io_ddr_out_ready),
    .io_ddr_out_valid(Scatters_15_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Scatters_15_io_ddr_out_bits_tdata),
    .io_end(Scatters_15_io_end)
  );
  Gather Gathers ( // @[nf_arm_doce_top_main.scala 37:23]
    .clock(Gathers_clock),
    .reset(Gathers_reset),
    .io_ddr_in_ready(Gathers_io_ddr_in_ready),
    .io_ddr_in_valid(Gathers_io_ddr_in_valid),
    .io_ddr_in_bits_tdata(Gathers_io_ddr_in_bits_tdata),
    .io_ddr_in_bits_tkeep(Gathers_io_ddr_in_bits_tkeep),
    .io_gather_out_0_ready(Gathers_io_gather_out_0_ready),
    .io_gather_out_0_valid(Gathers_io_gather_out_0_valid),
    .io_gather_out_0_bits_tdata(Gathers_io_gather_out_0_bits_tdata),
    .io_gather_out_1_ready(Gathers_io_gather_out_1_ready),
    .io_gather_out_1_valid(Gathers_io_gather_out_1_valid),
    .io_gather_out_1_bits_tdata(Gathers_io_gather_out_1_bits_tdata),
    .io_gather_out_2_ready(Gathers_io_gather_out_2_ready),
    .io_gather_out_2_valid(Gathers_io_gather_out_2_valid),
    .io_gather_out_2_bits_tdata(Gathers_io_gather_out_2_bits_tdata),
    .io_gather_out_3_ready(Gathers_io_gather_out_3_ready),
    .io_gather_out_3_valid(Gathers_io_gather_out_3_valid),
    .io_gather_out_3_bits_tdata(Gathers_io_gather_out_3_bits_tdata),
    .io_gather_out_4_ready(Gathers_io_gather_out_4_ready),
    .io_gather_out_4_valid(Gathers_io_gather_out_4_valid),
    .io_gather_out_4_bits_tdata(Gathers_io_gather_out_4_bits_tdata)
  );
  Apply Applys ( // @[nf_arm_doce_top_main.scala 38:22]
    .clock(Applys_clock),
    .reset(Applys_reset),
    .io_ddr_aw_ready(Applys_io_ddr_aw_ready),
    .io_ddr_aw_valid(Applys_io_ddr_aw_valid),
    .io_ddr_aw_bits_awaddr(Applys_io_ddr_aw_bits_awaddr),
    .io_ddr_aw_bits_awid(Applys_io_ddr_aw_bits_awid),
    .io_ddr_w_ready(Applys_io_ddr_w_ready),
    .io_ddr_w_valid(Applys_io_ddr_w_valid),
    .io_ddr_w_bits_wdata(Applys_io_ddr_w_bits_wdata),
    .io_ddr_w_bits_wstrb(Applys_io_ddr_w_bits_wstrb),
    .io_gather_in_ready(Applys_io_gather_in_ready),
    .io_gather_in_valid(Applys_io_gather_in_valid),
    .io_gather_in_bits_tdata(Applys_io_gather_in_bits_tdata),
    .io_level(Applys_io_level),
    .io_level_base_addr(Applys_io_level_base_addr),
    .io_end(Applys_io_end),
    .io_flush(Applys_io_flush)
  );
  Broadcast Broadcasts_0 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Broadcasts_0_clock),
    .reset(Broadcasts_0_reset),
    .io_ddr_ar_ready(Broadcasts_0_io_ddr_ar_ready),
    .io_ddr_ar_valid(Broadcasts_0_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Broadcasts_0_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Broadcasts_0_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Broadcasts_0_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Broadcasts_0_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Broadcasts_0_io_ddr_r_ready),
    .io_ddr_r_valid(Broadcasts_0_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Broadcasts_0_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Broadcasts_0_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Broadcasts_0_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Broadcasts_0_io_gather_in_ready),
    .io_gather_in_valid(Broadcasts_0_io_gather_in_valid),
    .io_gather_in_bits_tdata(Broadcasts_0_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Broadcasts_0_io_xbar_out_ready),
    .io_xbar_out_valid(Broadcasts_0_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Broadcasts_0_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Broadcasts_0_io_xbar_out_bits_tkeep),
    .io_embedding_base_addr(Broadcasts_0_io_embedding_base_addr),
    .io_edge_base_addr(Broadcasts_0_io_edge_base_addr),
    .io_signal(Broadcasts_0_io_signal),
    .io_traveled_edges(Broadcasts_0_io_traveled_edges),
    .io_start(Broadcasts_0_io_start),
    .io_root(Broadcasts_0_io_root),
    .io_issue_sync(Broadcasts_0_io_issue_sync),
    .io_recv_sync(Broadcasts_0_io_recv_sync)
  );
  Broadcast_1 Broadcasts_1 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Broadcasts_1_clock),
    .reset(Broadcasts_1_reset),
    .io_ddr_ar_ready(Broadcasts_1_io_ddr_ar_ready),
    .io_ddr_ar_valid(Broadcasts_1_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Broadcasts_1_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Broadcasts_1_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Broadcasts_1_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Broadcasts_1_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Broadcasts_1_io_ddr_r_ready),
    .io_ddr_r_valid(Broadcasts_1_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Broadcasts_1_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Broadcasts_1_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Broadcasts_1_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Broadcasts_1_io_gather_in_ready),
    .io_gather_in_valid(Broadcasts_1_io_gather_in_valid),
    .io_gather_in_bits_tdata(Broadcasts_1_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Broadcasts_1_io_xbar_out_ready),
    .io_xbar_out_valid(Broadcasts_1_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Broadcasts_1_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Broadcasts_1_io_xbar_out_bits_tkeep),
    .io_embedding_base_addr(Broadcasts_1_io_embedding_base_addr),
    .io_edge_base_addr(Broadcasts_1_io_edge_base_addr),
    .io_signal(Broadcasts_1_io_signal),
    .io_traveled_edges(Broadcasts_1_io_traveled_edges),
    .io_issue_sync(Broadcasts_1_io_issue_sync),
    .io_recv_sync(Broadcasts_1_io_recv_sync)
  );
  Broadcast_2 Broadcasts_2 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Broadcasts_2_clock),
    .reset(Broadcasts_2_reset),
    .io_ddr_ar_ready(Broadcasts_2_io_ddr_ar_ready),
    .io_ddr_ar_valid(Broadcasts_2_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Broadcasts_2_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Broadcasts_2_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Broadcasts_2_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Broadcasts_2_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Broadcasts_2_io_ddr_r_ready),
    .io_ddr_r_valid(Broadcasts_2_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Broadcasts_2_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Broadcasts_2_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Broadcasts_2_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Broadcasts_2_io_gather_in_ready),
    .io_gather_in_valid(Broadcasts_2_io_gather_in_valid),
    .io_gather_in_bits_tdata(Broadcasts_2_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Broadcasts_2_io_xbar_out_ready),
    .io_xbar_out_valid(Broadcasts_2_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Broadcasts_2_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Broadcasts_2_io_xbar_out_bits_tkeep),
    .io_embedding_base_addr(Broadcasts_2_io_embedding_base_addr),
    .io_edge_base_addr(Broadcasts_2_io_edge_base_addr),
    .io_signal(Broadcasts_2_io_signal),
    .io_traveled_edges(Broadcasts_2_io_traveled_edges),
    .io_issue_sync(Broadcasts_2_io_issue_sync),
    .io_recv_sync(Broadcasts_2_io_recv_sync)
  );
  Broadcast_3 Broadcasts_3 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Broadcasts_3_clock),
    .reset(Broadcasts_3_reset),
    .io_ddr_ar_ready(Broadcasts_3_io_ddr_ar_ready),
    .io_ddr_ar_valid(Broadcasts_3_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Broadcasts_3_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Broadcasts_3_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Broadcasts_3_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Broadcasts_3_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Broadcasts_3_io_ddr_r_ready),
    .io_ddr_r_valid(Broadcasts_3_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Broadcasts_3_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Broadcasts_3_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Broadcasts_3_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Broadcasts_3_io_gather_in_ready),
    .io_gather_in_valid(Broadcasts_3_io_gather_in_valid),
    .io_gather_in_bits_tdata(Broadcasts_3_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Broadcasts_3_io_xbar_out_ready),
    .io_xbar_out_valid(Broadcasts_3_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Broadcasts_3_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Broadcasts_3_io_xbar_out_bits_tkeep),
    .io_embedding_base_addr(Broadcasts_3_io_embedding_base_addr),
    .io_edge_base_addr(Broadcasts_3_io_edge_base_addr),
    .io_signal(Broadcasts_3_io_signal),
    .io_traveled_edges(Broadcasts_3_io_traveled_edges),
    .io_issue_sync(Broadcasts_3_io_issue_sync),
    .io_recv_sync(Broadcasts_3_io_recv_sync)
  );
  broadcast_xbar bxbar ( // @[nf_arm_doce_top_main.scala 43:21]
    .clock(bxbar_clock),
    .reset(bxbar_reset),
    .io_ddr_in_0_ready(bxbar_io_ddr_in_0_ready),
    .io_ddr_in_0_valid(bxbar_io_ddr_in_0_valid),
    .io_ddr_in_0_bits_tdata(bxbar_io_ddr_in_0_bits_tdata),
    .io_ddr_in_0_bits_tkeep(bxbar_io_ddr_in_0_bits_tkeep),
    .io_ddr_in_1_ready(bxbar_io_ddr_in_1_ready),
    .io_ddr_in_1_valid(bxbar_io_ddr_in_1_valid),
    .io_ddr_in_1_bits_tdata(bxbar_io_ddr_in_1_bits_tdata),
    .io_ddr_in_1_bits_tkeep(bxbar_io_ddr_in_1_bits_tkeep),
    .io_ddr_in_2_ready(bxbar_io_ddr_in_2_ready),
    .io_ddr_in_2_valid(bxbar_io_ddr_in_2_valid),
    .io_ddr_in_2_bits_tdata(bxbar_io_ddr_in_2_bits_tdata),
    .io_ddr_in_2_bits_tkeep(bxbar_io_ddr_in_2_bits_tkeep),
    .io_ddr_in_3_ready(bxbar_io_ddr_in_3_ready),
    .io_ddr_in_3_valid(bxbar_io_ddr_in_3_valid),
    .io_ddr_in_3_bits_tdata(bxbar_io_ddr_in_3_bits_tdata),
    .io_ddr_in_3_bits_tkeep(bxbar_io_ddr_in_3_bits_tkeep),
    .io_pe_out_0_ready(bxbar_io_pe_out_0_ready),
    .io_pe_out_0_valid(bxbar_io_pe_out_0_valid),
    .io_pe_out_0_bits_tdata(bxbar_io_pe_out_0_bits_tdata),
    .io_pe_out_0_bits_tkeep(bxbar_io_pe_out_0_bits_tkeep),
    .io_pe_out_1_ready(bxbar_io_pe_out_1_ready),
    .io_pe_out_1_valid(bxbar_io_pe_out_1_valid),
    .io_pe_out_1_bits_tdata(bxbar_io_pe_out_1_bits_tdata),
    .io_pe_out_1_bits_tkeep(bxbar_io_pe_out_1_bits_tkeep),
    .io_pe_out_2_ready(bxbar_io_pe_out_2_ready),
    .io_pe_out_2_valid(bxbar_io_pe_out_2_valid),
    .io_pe_out_2_bits_tdata(bxbar_io_pe_out_2_bits_tdata),
    .io_pe_out_2_bits_tkeep(bxbar_io_pe_out_2_bits_tkeep),
    .io_pe_out_3_ready(bxbar_io_pe_out_3_ready),
    .io_pe_out_3_valid(bxbar_io_pe_out_3_valid),
    .io_pe_out_3_bits_tdata(bxbar_io_pe_out_3_bits_tdata),
    .io_pe_out_3_bits_tkeep(bxbar_io_pe_out_3_bits_tkeep),
    .io_pe_out_4_ready(bxbar_io_pe_out_4_ready),
    .io_pe_out_4_valid(bxbar_io_pe_out_4_valid),
    .io_pe_out_4_bits_tdata(bxbar_io_pe_out_4_bits_tdata),
    .io_pe_out_4_bits_tkeep(bxbar_io_pe_out_4_bits_tkeep),
    .io_pe_out_5_ready(bxbar_io_pe_out_5_ready),
    .io_pe_out_5_valid(bxbar_io_pe_out_5_valid),
    .io_pe_out_5_bits_tdata(bxbar_io_pe_out_5_bits_tdata),
    .io_pe_out_5_bits_tkeep(bxbar_io_pe_out_5_bits_tkeep),
    .io_pe_out_6_ready(bxbar_io_pe_out_6_ready),
    .io_pe_out_6_valid(bxbar_io_pe_out_6_valid),
    .io_pe_out_6_bits_tdata(bxbar_io_pe_out_6_bits_tdata),
    .io_pe_out_6_bits_tkeep(bxbar_io_pe_out_6_bits_tkeep),
    .io_pe_out_7_ready(bxbar_io_pe_out_7_ready),
    .io_pe_out_7_valid(bxbar_io_pe_out_7_valid),
    .io_pe_out_7_bits_tdata(bxbar_io_pe_out_7_bits_tdata),
    .io_pe_out_7_bits_tkeep(bxbar_io_pe_out_7_bits_tkeep),
    .io_pe_out_8_ready(bxbar_io_pe_out_8_ready),
    .io_pe_out_8_valid(bxbar_io_pe_out_8_valid),
    .io_pe_out_8_bits_tdata(bxbar_io_pe_out_8_bits_tdata),
    .io_pe_out_8_bits_tkeep(bxbar_io_pe_out_8_bits_tkeep),
    .io_pe_out_9_ready(bxbar_io_pe_out_9_ready),
    .io_pe_out_9_valid(bxbar_io_pe_out_9_valid),
    .io_pe_out_9_bits_tdata(bxbar_io_pe_out_9_bits_tdata),
    .io_pe_out_9_bits_tkeep(bxbar_io_pe_out_9_bits_tkeep),
    .io_pe_out_10_ready(bxbar_io_pe_out_10_ready),
    .io_pe_out_10_valid(bxbar_io_pe_out_10_valid),
    .io_pe_out_10_bits_tdata(bxbar_io_pe_out_10_bits_tdata),
    .io_pe_out_10_bits_tkeep(bxbar_io_pe_out_10_bits_tkeep),
    .io_pe_out_11_ready(bxbar_io_pe_out_11_ready),
    .io_pe_out_11_valid(bxbar_io_pe_out_11_valid),
    .io_pe_out_11_bits_tdata(bxbar_io_pe_out_11_bits_tdata),
    .io_pe_out_11_bits_tkeep(bxbar_io_pe_out_11_bits_tkeep),
    .io_pe_out_12_ready(bxbar_io_pe_out_12_ready),
    .io_pe_out_12_valid(bxbar_io_pe_out_12_valid),
    .io_pe_out_12_bits_tdata(bxbar_io_pe_out_12_bits_tdata),
    .io_pe_out_12_bits_tkeep(bxbar_io_pe_out_12_bits_tkeep),
    .io_pe_out_13_ready(bxbar_io_pe_out_13_ready),
    .io_pe_out_13_valid(bxbar_io_pe_out_13_valid),
    .io_pe_out_13_bits_tdata(bxbar_io_pe_out_13_bits_tdata),
    .io_pe_out_13_bits_tkeep(bxbar_io_pe_out_13_bits_tkeep),
    .io_pe_out_14_ready(bxbar_io_pe_out_14_ready),
    .io_pe_out_14_valid(bxbar_io_pe_out_14_valid),
    .io_pe_out_14_bits_tdata(bxbar_io_pe_out_14_bits_tdata),
    .io_pe_out_14_bits_tkeep(bxbar_io_pe_out_14_bits_tkeep),
    .io_pe_out_15_ready(bxbar_io_pe_out_15_ready),
    .io_pe_out_15_valid(bxbar_io_pe_out_15_valid),
    .io_pe_out_15_bits_tdata(bxbar_io_pe_out_15_bits_tdata),
    .io_pe_out_15_bits_tkeep(bxbar_io_pe_out_15_bits_tkeep)
  );
  assign io_config_awready = controls_io_config_awready; // @[nf_arm_doce_top_main.scala 90:22]
  assign io_config_arready = controls_io_config_arready; // @[nf_arm_doce_top_main.scala 90:22]
  assign io_config_wready = controls_io_config_wready; // @[nf_arm_doce_top_main.scala 90:22]
  assign io_config_rdata = controls_io_config_rdata; // @[nf_arm_doce_top_main.scala 90:22]
  assign io_config_rresp = 2'h0; // @[nf_arm_doce_top_main.scala 90:22]
  assign io_config_rvalid = controls_io_config_rvalid; // @[nf_arm_doce_top_main.scala 90:22]
  assign io_config_bresp = 2'h0; // @[nf_arm_doce_top_main.scala 90:22]
  assign io_config_bvalid = controls_io_config_bvalid; // @[nf_arm_doce_top_main.scala 90:22]
  assign io_PLmemory_0_aw_valid = pl_mc_io_ddr_out_0_aw_valid; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_aw_bits_awaddr = pl_mc_io_ddr_out_0_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_aw_bits_awid = 7'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_aw_bits_awlen = 8'hf; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_aw_bits_awsize = 3'h6; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_ar_valid = pl_mc_io_ddr_out_0_ar_valid; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_ar_bits_araddr = pl_mc_io_ddr_out_0_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_ar_bits_arid = 7'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_ar_bits_arlen = 8'hf; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_ar_bits_arsize = 3'h6; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_w_valid = pl_mc_io_ddr_out_0_w_valid; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_w_bits_wdata = pl_mc_io_ddr_out_0_w_bits_wdata; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_w_bits_wstrb = 64'hffffffffffffffff; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_w_bits_wlast = pl_mc_io_ddr_out_0_w_bits_wlast; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_r_ready = 1'h1; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_0_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_aw_valid = pl_mc_io_ddr_out_1_aw_valid; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_aw_bits_awaddr = pl_mc_io_ddr_out_1_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_aw_bits_awid = pl_mc_io_ddr_out_1_aw_bits_awid; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_aw_bits_awsize = 3'h2; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_ar_valid = 1'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_ar_bits_araddr = 64'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_ar_bits_arid = 7'h40; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_ar_bits_arlen = 8'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_ar_bits_arsize = 3'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_ar_bits_arburst = 2'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_w_valid = pl_mc_io_ddr_out_1_w_valid; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_w_bits_wdata = pl_mc_io_ddr_out_1_w_bits_wdata; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_w_bits_wstrb = pl_mc_io_ddr_out_1_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_w_bits_wlast = 1'h1; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_r_ready = 1'h0; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PLmemory_1_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 45:15]
  assign io_PSmemory_0_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 75:18]
  assign io_PSmemory_0_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 46:12]
  assign io_PSmemory_0_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 47:10]
  assign io_PSmemory_0_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 48:11]
  assign io_PSmemory_0_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 49:12]
  assign io_PSmemory_0_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 50:13]
  assign io_PSmemory_0_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_0_ar_valid = Broadcasts_0_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_0_ar_bits_araddr = Broadcasts_0_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_0_ar_bits_arid = Broadcasts_0_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_0_ar_bits_arlen = Broadcasts_0_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_0_ar_bits_arsize = Broadcasts_0_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_0_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_0_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_0_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 77:17]
  assign io_PSmemory_0_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 61:11]
  assign io_PSmemory_0_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 62:11]
  assign io_PSmemory_0_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 63:11]
  assign io_PSmemory_0_r_ready = Broadcasts_0_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 56:18]
  assign io_PSmemory_0_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 73:17]
  assign io_PSmemory_1_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 75:18]
  assign io_PSmemory_1_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 46:12]
  assign io_PSmemory_1_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 47:10]
  assign io_PSmemory_1_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 48:11]
  assign io_PSmemory_1_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 49:12]
  assign io_PSmemory_1_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 50:13]
  assign io_PSmemory_1_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_1_ar_valid = Broadcasts_1_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_1_ar_bits_araddr = Broadcasts_1_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_1_ar_bits_arid = Broadcasts_1_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_1_ar_bits_arlen = Broadcasts_1_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_1_ar_bits_arsize = Broadcasts_1_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_1_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_1_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_1_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 77:17]
  assign io_PSmemory_1_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 61:11]
  assign io_PSmemory_1_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 62:11]
  assign io_PSmemory_1_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 63:11]
  assign io_PSmemory_1_r_ready = Broadcasts_1_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 56:18]
  assign io_PSmemory_1_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 73:17]
  assign io_PSmemory_2_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 75:18]
  assign io_PSmemory_2_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 46:12]
  assign io_PSmemory_2_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 47:10]
  assign io_PSmemory_2_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 48:11]
  assign io_PSmemory_2_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 49:12]
  assign io_PSmemory_2_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 50:13]
  assign io_PSmemory_2_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_2_ar_valid = Broadcasts_2_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_2_ar_bits_araddr = Broadcasts_2_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_2_ar_bits_arid = Broadcasts_2_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_2_ar_bits_arlen = Broadcasts_2_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_2_ar_bits_arsize = Broadcasts_2_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_2_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_2_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_2_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 77:17]
  assign io_PSmemory_2_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 61:11]
  assign io_PSmemory_2_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 62:11]
  assign io_PSmemory_2_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 63:11]
  assign io_PSmemory_2_r_ready = Broadcasts_2_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 56:18]
  assign io_PSmemory_2_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 73:17]
  assign io_PSmemory_3_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 75:18]
  assign io_PSmemory_3_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 46:12]
  assign io_PSmemory_3_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 47:10]
  assign io_PSmemory_3_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 48:11]
  assign io_PSmemory_3_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 49:12]
  assign io_PSmemory_3_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 50:13]
  assign io_PSmemory_3_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_3_ar_valid = Broadcasts_3_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_3_ar_bits_araddr = Broadcasts_3_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_3_ar_bits_arid = Broadcasts_3_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_3_ar_bits_arlen = Broadcasts_3_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_3_ar_bits_arsize = Broadcasts_3_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_3_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_3_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 57:19]
  assign io_PSmemory_3_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 77:17]
  assign io_PSmemory_3_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 61:11]
  assign io_PSmemory_3_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 62:11]
  assign io_PSmemory_3_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 63:11]
  assign io_PSmemory_3_r_ready = Broadcasts_3_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 56:18]
  assign io_PSmemory_3_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 73:17]
  assign controls_clock = clock;
  assign controls_reset = reset;
  assign controls_io_fin_0 = Scatters_0_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_1 = Scatters_1_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_2 = Scatters_2_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_3 = Scatters_3_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_4 = Scatters_4_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_5 = Scatters_5_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_6 = Scatters_6_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_7 = Scatters_7_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_8 = Scatters_8_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_9 = Scatters_9_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_10 = Scatters_10_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_11 = Scatters_11_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_12 = Scatters_12_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_13 = Scatters_13_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_14 = Scatters_14_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_fin_15 = Scatters_15_io_end; // @[nf_arm_doce_top_main.scala 66:26]
  assign controls_io_unvisited_size = pl_mc_io_unvisited_size; // @[nf_arm_doce_top_main.scala 92:30]
  assign controls_io_traveled_edges = _controls_io_traveled_edges_T_3 + Broadcasts_3_io_traveled_edges; // @[nf_arm_doce_top_main.scala 91:82]
  assign controls_io_config_awaddr = io_config_awaddr; // @[nf_arm_doce_top_main.scala 90:22]
  assign controls_io_config_araddr = io_config_araddr; // @[nf_arm_doce_top_main.scala 90:22]
  assign controls_io_config_arvalid = io_config_arvalid; // @[nf_arm_doce_top_main.scala 90:22]
  assign controls_io_config_wdata = io_config_wdata; // @[nf_arm_doce_top_main.scala 90:22]
  assign controls_io_config_wstrb = io_config_wstrb; // @[nf_arm_doce_top_main.scala 90:22]
  assign controls_io_config_wvalid = io_config_wvalid; // @[nf_arm_doce_top_main.scala 90:22]
  assign controls_io_config_rready = io_config_rready; // @[nf_arm_doce_top_main.scala 90:22]
  assign controls_io_config_bready = io_config_bready; // @[nf_arm_doce_top_main.scala 90:22]
  assign controls_io_flush_cache_end = Applys_io_end; // @[nf_arm_doce_top_main.scala 93:31]
  assign pl_mc_clock = clock;
  assign pl_mc_reset = reset;
  assign pl_mc_io_cacheable_out_ready = Gathers_io_ddr_in_ready; // @[nf_arm_doce_top_main.scala 46:21]
  assign pl_mc_io_cacheable_in_0_valid = Scatters_0_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_0_bits_tdata = Scatters_0_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_1_valid = Scatters_1_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_1_bits_tdata = Scatters_1_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_2_valid = Scatters_2_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_2_bits_tdata = Scatters_2_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_3_valid = Scatters_3_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_3_bits_tdata = Scatters_3_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_4_valid = Scatters_4_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_4_bits_tdata = Scatters_4_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_5_valid = Scatters_5_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_5_bits_tdata = Scatters_5_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_6_valid = Scatters_6_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_6_bits_tdata = Scatters_6_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_7_valid = Scatters_7_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_7_bits_tdata = Scatters_7_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_8_valid = Scatters_8_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_8_bits_tdata = Scatters_8_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_9_valid = Scatters_9_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_9_bits_tdata = Scatters_9_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_10_valid = Scatters_10_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_10_bits_tdata = Scatters_10_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_11_valid = Scatters_11_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_11_bits_tdata = Scatters_11_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_12_valid = Scatters_12_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_12_bits_tdata = Scatters_12_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_13_valid = Scatters_13_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_13_bits_tdata = Scatters_13_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_14_valid = Scatters_14_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_14_bits_tdata = Scatters_14_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_15_valid = Scatters_15_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_cacheable_in_15_bits_tdata = Scatters_15_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:21]
  assign pl_mc_io_non_cacheable_in_aw_valid = Applys_io_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 50:20]
  assign pl_mc_io_non_cacheable_in_aw_bits_awaddr = Applys_io_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 50:20]
  assign pl_mc_io_non_cacheable_in_aw_bits_awid = Applys_io_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 50:20]
  assign pl_mc_io_non_cacheable_in_w_valid = Applys_io_ddr_w_valid; // @[nf_arm_doce_top_main.scala 49:19]
  assign pl_mc_io_non_cacheable_in_w_bits_wdata = Applys_io_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 49:19]
  assign pl_mc_io_non_cacheable_in_w_bits_wstrb = Applys_io_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 49:19]
  assign pl_mc_io_ddr_out_0_aw_ready = io_PLmemory_0_aw_ready; // @[nf_arm_doce_top_main.scala 45:15]
  assign pl_mc_io_ddr_out_0_ar_ready = io_PLmemory_0_ar_ready; // @[nf_arm_doce_top_main.scala 45:15]
  assign pl_mc_io_ddr_out_0_w_ready = io_PLmemory_0_w_ready; // @[nf_arm_doce_top_main.scala 45:15]
  assign pl_mc_io_ddr_out_0_r_valid = io_PLmemory_0_r_valid; // @[nf_arm_doce_top_main.scala 45:15]
  assign pl_mc_io_ddr_out_0_r_bits_rdata = io_PLmemory_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 45:15]
  assign pl_mc_io_ddr_out_0_r_bits_rlast = io_PLmemory_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 45:15]
  assign pl_mc_io_ddr_out_1_aw_ready = io_PLmemory_1_aw_ready; // @[nf_arm_doce_top_main.scala 45:15]
  assign pl_mc_io_ddr_out_1_w_ready = io_PLmemory_1_w_ready; // @[nf_arm_doce_top_main.scala 45:15]
  assign pl_mc_io_tiers_base_addr_0 = {controls_io_data_9,controls_io_data_8}; // @[Cat.scala 30:58]
  assign pl_mc_io_tiers_base_addr_1 = {controls_io_data_11,controls_io_data_10}; // @[Cat.scala 30:58]
  assign pl_mc_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 114:18]
  assign pl_mc_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 113:19]
  assign pl_mc_io_end = controls_io_data_0[1]; // @[nf_arm_doce_top_main.scala 115:38]
  assign Scatters_0_clock = clock;
  assign Scatters_0_reset = reset;
  assign Scatters_0_io_xbar_in_valid = bxbar_io_pe_out_0_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_0_io_xbar_in_bits_tdata = bxbar_io_pe_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_0_io_xbar_in_bits_tkeep = bxbar_io_pe_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_0_io_ddr_out_ready = pl_mc_io_cacheable_in_0_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_1_clock = clock;
  assign Scatters_1_reset = reset;
  assign Scatters_1_io_xbar_in_valid = bxbar_io_pe_out_1_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_1_io_xbar_in_bits_tdata = bxbar_io_pe_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_1_io_xbar_in_bits_tkeep = bxbar_io_pe_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_1_io_ddr_out_ready = pl_mc_io_cacheable_in_1_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_2_clock = clock;
  assign Scatters_2_reset = reset;
  assign Scatters_2_io_xbar_in_valid = bxbar_io_pe_out_2_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_2_io_xbar_in_bits_tdata = bxbar_io_pe_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_2_io_xbar_in_bits_tkeep = bxbar_io_pe_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_2_io_ddr_out_ready = pl_mc_io_cacheable_in_2_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_3_clock = clock;
  assign Scatters_3_reset = reset;
  assign Scatters_3_io_xbar_in_valid = bxbar_io_pe_out_3_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_3_io_xbar_in_bits_tdata = bxbar_io_pe_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_3_io_xbar_in_bits_tkeep = bxbar_io_pe_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_3_io_ddr_out_ready = pl_mc_io_cacheable_in_3_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_4_clock = clock;
  assign Scatters_4_reset = reset;
  assign Scatters_4_io_xbar_in_valid = bxbar_io_pe_out_4_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_4_io_xbar_in_bits_tdata = bxbar_io_pe_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_4_io_xbar_in_bits_tkeep = bxbar_io_pe_out_4_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_4_io_ddr_out_ready = pl_mc_io_cacheable_in_4_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_5_clock = clock;
  assign Scatters_5_reset = reset;
  assign Scatters_5_io_xbar_in_valid = bxbar_io_pe_out_5_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_5_io_xbar_in_bits_tdata = bxbar_io_pe_out_5_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_5_io_xbar_in_bits_tkeep = bxbar_io_pe_out_5_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_5_io_ddr_out_ready = pl_mc_io_cacheable_in_5_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_6_clock = clock;
  assign Scatters_6_reset = reset;
  assign Scatters_6_io_xbar_in_valid = bxbar_io_pe_out_6_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_6_io_xbar_in_bits_tdata = bxbar_io_pe_out_6_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_6_io_xbar_in_bits_tkeep = bxbar_io_pe_out_6_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_6_io_ddr_out_ready = pl_mc_io_cacheable_in_6_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_7_clock = clock;
  assign Scatters_7_reset = reset;
  assign Scatters_7_io_xbar_in_valid = bxbar_io_pe_out_7_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_7_io_xbar_in_bits_tdata = bxbar_io_pe_out_7_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_7_io_xbar_in_bits_tkeep = bxbar_io_pe_out_7_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_7_io_ddr_out_ready = pl_mc_io_cacheable_in_7_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_8_clock = clock;
  assign Scatters_8_reset = reset;
  assign Scatters_8_io_xbar_in_valid = bxbar_io_pe_out_8_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_8_io_xbar_in_bits_tdata = bxbar_io_pe_out_8_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_8_io_xbar_in_bits_tkeep = bxbar_io_pe_out_8_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_8_io_ddr_out_ready = pl_mc_io_cacheable_in_8_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_9_clock = clock;
  assign Scatters_9_reset = reset;
  assign Scatters_9_io_xbar_in_valid = bxbar_io_pe_out_9_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_9_io_xbar_in_bits_tdata = bxbar_io_pe_out_9_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_9_io_xbar_in_bits_tkeep = bxbar_io_pe_out_9_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_9_io_ddr_out_ready = pl_mc_io_cacheable_in_9_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_10_clock = clock;
  assign Scatters_10_reset = reset;
  assign Scatters_10_io_xbar_in_valid = bxbar_io_pe_out_10_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_10_io_xbar_in_bits_tdata = bxbar_io_pe_out_10_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_10_io_xbar_in_bits_tkeep = bxbar_io_pe_out_10_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_10_io_ddr_out_ready = pl_mc_io_cacheable_in_10_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_11_clock = clock;
  assign Scatters_11_reset = reset;
  assign Scatters_11_io_xbar_in_valid = bxbar_io_pe_out_11_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_11_io_xbar_in_bits_tdata = bxbar_io_pe_out_11_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_11_io_xbar_in_bits_tkeep = bxbar_io_pe_out_11_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_11_io_ddr_out_ready = pl_mc_io_cacheable_in_11_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_12_clock = clock;
  assign Scatters_12_reset = reset;
  assign Scatters_12_io_xbar_in_valid = bxbar_io_pe_out_12_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_12_io_xbar_in_bits_tdata = bxbar_io_pe_out_12_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_12_io_xbar_in_bits_tkeep = bxbar_io_pe_out_12_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_12_io_ddr_out_ready = pl_mc_io_cacheable_in_12_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_13_clock = clock;
  assign Scatters_13_reset = reset;
  assign Scatters_13_io_xbar_in_valid = bxbar_io_pe_out_13_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_13_io_xbar_in_bits_tdata = bxbar_io_pe_out_13_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_13_io_xbar_in_bits_tkeep = bxbar_io_pe_out_13_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_13_io_ddr_out_ready = pl_mc_io_cacheable_in_13_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_14_clock = clock;
  assign Scatters_14_reset = reset;
  assign Scatters_14_io_xbar_in_valid = bxbar_io_pe_out_14_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_14_io_xbar_in_bits_tdata = bxbar_io_pe_out_14_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_14_io_xbar_in_bits_tkeep = bxbar_io_pe_out_14_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_14_io_ddr_out_ready = pl_mc_io_cacheable_in_14_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Scatters_15_clock = clock;
  assign Scatters_15_reset = reset;
  assign Scatters_15_io_xbar_in_valid = bxbar_io_pe_out_15_valid; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_15_io_xbar_in_bits_tdata = bxbar_io_pe_out_15_bits_tdata; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_15_io_xbar_in_bits_tkeep = bxbar_io_pe_out_15_bits_tkeep; // @[nf_arm_doce_top_main.scala 64:21]
  assign Scatters_15_io_ddr_out_ready = pl_mc_io_cacheable_in_15_ready; // @[nf_arm_doce_top_main.scala 65:21]
  assign Gathers_clock = clock;
  assign Gathers_reset = reset;
  assign Gathers_io_ddr_in_valid = pl_mc_io_cacheable_out_valid; // @[nf_arm_doce_top_main.scala 46:21]
  assign Gathers_io_ddr_in_bits_tdata = pl_mc_io_cacheable_out_bits_tdata; // @[nf_arm_doce_top_main.scala 46:21]
  assign Gathers_io_ddr_in_bits_tkeep = pl_mc_io_cacheable_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 46:21]
  assign Gathers_io_gather_out_0_ready = Broadcasts_0_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 55:22]
  assign Gathers_io_gather_out_1_ready = Broadcasts_1_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 55:22]
  assign Gathers_io_gather_out_2_ready = Broadcasts_2_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 55:22]
  assign Gathers_io_gather_out_3_ready = Broadcasts_3_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 55:22]
  assign Gathers_io_gather_out_4_ready = Applys_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 48:23]
  assign Applys_clock = clock;
  assign Applys_reset = reset;
  assign Applys_io_ddr_aw_ready = pl_mc_io_non_cacheable_in_aw_ready; // @[nf_arm_doce_top_main.scala 50:20]
  assign Applys_io_ddr_w_ready = pl_mc_io_non_cacheable_in_w_ready; // @[nf_arm_doce_top_main.scala 49:19]
  assign Applys_io_gather_in_valid = Gathers_io_gather_out_4_valid; // @[nf_arm_doce_top_main.scala 48:23]
  assign Applys_io_gather_in_bits_tdata = Gathers_io_gather_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 48:23]
  assign Applys_io_level = controls_io_level; // @[nf_arm_doce_top_main.scala 97:19]
  assign Applys_io_level_base_addr = {controls_io_data_6,controls_io_data_5}; // @[Cat.scala 30:58]
  assign Applys_io_flush = controls_io_flush_cache; // @[nf_arm_doce_top_main.scala 95:19]
  assign Broadcasts_0_clock = clock;
  assign Broadcasts_0_reset = reset;
  assign Broadcasts_0_io_ddr_ar_ready = io_PSmemory_0_ar_ready; // @[nf_arm_doce_top_main.scala 57:19]
  assign Broadcasts_0_io_ddr_r_valid = io_PSmemory_0_r_valid; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_0_io_ddr_r_bits_rdata = io_PSmemory_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_0_io_ddr_r_bits_rid = io_PSmemory_0_r_bits_rid; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_0_io_ddr_r_bits_rlast = io_PSmemory_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_0_io_gather_in_valid = Gathers_io_gather_out_0_valid; // @[nf_arm_doce_top_main.scala 55:22]
  assign Broadcasts_0_io_gather_in_bits_tdata = Gathers_io_gather_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 55:22]
  assign Broadcasts_0_io_xbar_out_ready = bxbar_io_ddr_in_0_ready; // @[nf_arm_doce_top_main.scala 58:26]
  assign Broadcasts_0_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Broadcasts_0_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Broadcasts_0_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 101:19]
  assign Broadcasts_0_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 105:20]
  assign Broadcasts_0_io_root = controls_io_data_7; // @[nf_arm_doce_top_main.scala 100:17]
  assign Broadcasts_0_io_recv_sync = {Broadcasts_0_io_recv_sync_hi,Broadcasts_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 59:77]
  assign Broadcasts_1_clock = clock;
  assign Broadcasts_1_reset = reset;
  assign Broadcasts_1_io_ddr_ar_ready = io_PSmemory_1_ar_ready; // @[nf_arm_doce_top_main.scala 57:19]
  assign Broadcasts_1_io_ddr_r_valid = io_PSmemory_1_r_valid; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_1_io_ddr_r_bits_rdata = io_PSmemory_1_r_bits_rdata; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_1_io_ddr_r_bits_rid = io_PSmemory_1_r_bits_rid; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_1_io_ddr_r_bits_rlast = io_PSmemory_1_r_bits_rlast; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_1_io_gather_in_valid = Gathers_io_gather_out_1_valid; // @[nf_arm_doce_top_main.scala 55:22]
  assign Broadcasts_1_io_gather_in_bits_tdata = Gathers_io_gather_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 55:22]
  assign Broadcasts_1_io_xbar_out_ready = bxbar_io_ddr_in_1_ready; // @[nf_arm_doce_top_main.scala 58:26]
  assign Broadcasts_1_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Broadcasts_1_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Broadcasts_1_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 101:19]
  assign Broadcasts_1_io_recv_sync = {Broadcasts_0_io_recv_sync_hi,Broadcasts_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 59:77]
  assign Broadcasts_2_clock = clock;
  assign Broadcasts_2_reset = reset;
  assign Broadcasts_2_io_ddr_ar_ready = io_PSmemory_2_ar_ready; // @[nf_arm_doce_top_main.scala 57:19]
  assign Broadcasts_2_io_ddr_r_valid = io_PSmemory_2_r_valid; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_2_io_ddr_r_bits_rdata = io_PSmemory_2_r_bits_rdata; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_2_io_ddr_r_bits_rid = io_PSmemory_2_r_bits_rid; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_2_io_ddr_r_bits_rlast = io_PSmemory_2_r_bits_rlast; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_2_io_gather_in_valid = Gathers_io_gather_out_2_valid; // @[nf_arm_doce_top_main.scala 55:22]
  assign Broadcasts_2_io_gather_in_bits_tdata = Gathers_io_gather_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 55:22]
  assign Broadcasts_2_io_xbar_out_ready = bxbar_io_ddr_in_2_ready; // @[nf_arm_doce_top_main.scala 58:26]
  assign Broadcasts_2_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Broadcasts_2_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Broadcasts_2_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 101:19]
  assign Broadcasts_2_io_recv_sync = {Broadcasts_0_io_recv_sync_hi,Broadcasts_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 59:77]
  assign Broadcasts_3_clock = clock;
  assign Broadcasts_3_reset = reset;
  assign Broadcasts_3_io_ddr_ar_ready = io_PSmemory_3_ar_ready; // @[nf_arm_doce_top_main.scala 57:19]
  assign Broadcasts_3_io_ddr_r_valid = io_PSmemory_3_r_valid; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_3_io_ddr_r_bits_rdata = io_PSmemory_3_r_bits_rdata; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_3_io_ddr_r_bits_rid = io_PSmemory_3_r_bits_rid; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_3_io_ddr_r_bits_rlast = io_PSmemory_3_r_bits_rlast; // @[nf_arm_doce_top_main.scala 56:18]
  assign Broadcasts_3_io_gather_in_valid = Gathers_io_gather_out_3_valid; // @[nf_arm_doce_top_main.scala 55:22]
  assign Broadcasts_3_io_gather_in_bits_tdata = Gathers_io_gather_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 55:22]
  assign Broadcasts_3_io_xbar_out_ready = bxbar_io_ddr_in_3_ready; // @[nf_arm_doce_top_main.scala 58:26]
  assign Broadcasts_3_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Broadcasts_3_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Broadcasts_3_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 101:19]
  assign Broadcasts_3_io_recv_sync = {Broadcasts_0_io_recv_sync_hi,Broadcasts_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 59:77]
  assign bxbar_clock = clock;
  assign bxbar_reset = reset;
  assign bxbar_io_ddr_in_0_valid = Broadcasts_0_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_0_bits_tdata = Broadcasts_0_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_0_bits_tkeep = Broadcasts_0_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_1_valid = Broadcasts_1_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_1_bits_tdata = Broadcasts_1_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_1_bits_tkeep = Broadcasts_1_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_2_valid = Broadcasts_2_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_2_bits_tdata = Broadcasts_2_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_2_bits_tkeep = Broadcasts_2_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_3_valid = Broadcasts_3_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_3_bits_tdata = Broadcasts_3_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_ddr_in_3_bits_tkeep = Broadcasts_3_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 58:26]
  assign bxbar_io_pe_out_0_ready = Scatters_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_1_ready = Scatters_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_2_ready = Scatters_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_3_ready = Scatters_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_4_ready = Scatters_4_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_5_ready = Scatters_5_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_6_ready = Scatters_6_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_7_ready = Scatters_7_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_8_ready = Scatters_8_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_9_ready = Scatters_9_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_10_ready = Scatters_10_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_11_ready = Scatters_11_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_12_ready = Scatters_12_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_13_ready = Scatters_13_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_14_ready = Scatters_14_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
  assign bxbar_io_pe_out_15_ready = Scatters_15_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 64:21]
endmodule
