module LookupTable(
  input         clock,
  input         reset,
  output [31:0] io_data_0,
  output [31:0] io_data_1,
  output [31:0] io_data_2,
  output [31:0] io_data_3,
  output [31:0] io_data_4,
  output [31:0] io_data_5,
  output [31:0] io_data_6,
  output [31:0] io_data_7,
  output [31:0] io_data_8,
  output [31:0] io_data_9,
  output [31:0] io_data_10,
  output [31:0] io_data_11,
  output [31:0] io_data_12,
  output [31:0] io_data_13,
  output [31:0] io_data_16,
  output [31:0] io_data_17,
  output [31:0] io_data_18,
  input  [31:0] io_dataIn_0,
  input  [31:0] io_dataIn_1,
  input         io_writeFlag_0,
  input         io_writeFlag_1,
  input  [4:0]  io_wptr_0,
  input  [4:0]  io_wptr_1,
  input  [63:0] config_awaddr,
  input         config_awvalid,
  output        config_awready,
  input  [63:0] config_araddr,
  input         config_arvalid,
  output        config_arready,
  input  [31:0] config_wdata,
  input         config_wvalid,
  output        config_wready,
  output [31:0] config_rdata,
  output        config_rvalid,
  input         config_rready,
  output        config_bvalid,
  input         config_bready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] table_0; // @[util.scala 16:22]
  reg [31:0] table_1; // @[util.scala 16:22]
  reg [31:0] table_2; // @[util.scala 16:22]
  reg [31:0] table_3; // @[util.scala 16:22]
  reg [31:0] table_4; // @[util.scala 16:22]
  reg [31:0] table_5; // @[util.scala 16:22]
  reg [31:0] table_6; // @[util.scala 16:22]
  reg [31:0] table_7; // @[util.scala 16:22]
  reg [31:0] table_8; // @[util.scala 16:22]
  reg [31:0] table_9; // @[util.scala 16:22]
  reg [31:0] table_10; // @[util.scala 16:22]
  reg [31:0] table_11; // @[util.scala 16:22]
  reg [31:0] table_12; // @[util.scala 16:22]
  reg [31:0] table_13; // @[util.scala 16:22]
  reg [31:0] table_14; // @[util.scala 16:22]
  reg [31:0] table_15; // @[util.scala 16:22]
  reg [31:0] table_16; // @[util.scala 16:22]
  reg [31:0] table_17; // @[util.scala 16:22]
  reg [31:0] table_18; // @[util.scala 16:22]
  reg [31:0] table_19; // @[util.scala 16:22]
  reg [31:0] table_20; // @[util.scala 16:22]
  reg [31:0] table_21; // @[util.scala 16:22]
  reg [31:0] table_22; // @[util.scala 16:22]
  reg [31:0] table_23; // @[util.scala 16:22]
  reg [31:0] table_24; // @[util.scala 16:22]
  reg [31:0] table_25; // @[util.scala 16:22]
  reg [31:0] table_26; // @[util.scala 16:22]
  reg [31:0] table_27; // @[util.scala 16:22]
  reg [31:0] table_28; // @[util.scala 16:22]
  reg [31:0] table_29; // @[util.scala 16:22]
  reg [31:0] table_30; // @[util.scala 16:22]
  reg [31:0] table_31; // @[util.scala 16:22]
  reg [2:0] status; // @[util.scala 26:23]
  wire [2:0] _GEN_3 = config_bready ? 3'h0 : status; // @[util.scala 41:24 util.scala 42:14 util.scala 26:23]
  wire [2:0] _GEN_4 = config_rready ? 3'h0 : status; // @[util.scala 47:25 util.scala 48:14 util.scala 26:23]
  wire [2:0] _GEN_5 = status == 3'h5 ? _GEN_4 : status; // @[util.scala 46:36 util.scala 26:23]
  wire [2:0] _GEN_6 = status == 3'h4 ? 3'h5 : _GEN_5; // @[util.scala 44:35 util.scala 45:12]
  wire [2:0] _GEN_7 = status == 3'h3 ? _GEN_3 : _GEN_6; // @[util.scala 40:35]
  wire  wvalid = config_wvalid & config_wready; // @[util.scala 64:30]
  reg [4:0] ewaddr; // @[util.scala 65:19]
  wire  _T_7 = io_writeFlag_0 & io_writeFlag_1; // @[util.scala 70:39]
  wire [31:0] _GEN_12 = 5'h0 == ewaddr ? config_wdata : table_0; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_13 = 5'h1 == ewaddr ? config_wdata : table_1; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_14 = 5'h2 == ewaddr ? config_wdata : table_2; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_15 = 5'h3 == ewaddr ? config_wdata : table_3; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_16 = 5'h4 == ewaddr ? config_wdata : table_4; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_17 = 5'h5 == ewaddr ? config_wdata : table_5; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_18 = 5'h6 == ewaddr ? config_wdata : table_6; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_19 = 5'h7 == ewaddr ? config_wdata : table_7; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_20 = 5'h8 == ewaddr ? config_wdata : table_8; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_21 = 5'h9 == ewaddr ? config_wdata : table_9; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_22 = 5'ha == ewaddr ? config_wdata : table_10; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_23 = 5'hb == ewaddr ? config_wdata : table_11; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_24 = 5'hc == ewaddr ? config_wdata : table_12; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_25 = 5'hd == ewaddr ? config_wdata : table_13; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_26 = 5'he == ewaddr ? config_wdata : table_14; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_27 = 5'hf == ewaddr ? config_wdata : table_15; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_28 = 5'h10 == ewaddr ? config_wdata : table_16; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_29 = 5'h11 == ewaddr ? config_wdata : table_17; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_30 = 5'h12 == ewaddr ? config_wdata : table_18; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_31 = 5'h13 == ewaddr ? config_wdata : table_19; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_32 = 5'h14 == ewaddr ? config_wdata : table_20; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_33 = 5'h15 == ewaddr ? config_wdata : table_21; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_34 = 5'h16 == ewaddr ? config_wdata : table_22; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_35 = 5'h17 == ewaddr ? config_wdata : table_23; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_36 = 5'h18 == ewaddr ? config_wdata : table_24; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_37 = 5'h19 == ewaddr ? config_wdata : table_25; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_38 = 5'h1a == ewaddr ? config_wdata : table_26; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_39 = 5'h1b == ewaddr ? config_wdata : table_27; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_40 = 5'h1c == ewaddr ? config_wdata : table_28; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_41 = 5'h1d == ewaddr ? config_wdata : table_29; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_42 = 5'h1e == ewaddr ? config_wdata : table_30; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_43 = 5'h1f == ewaddr ? config_wdata : table_31; // @[util.scala 71:19 util.scala 71:19 util.scala 16:22]
  wire [31:0] _GEN_44 = 5'h0 == io_wptr_0 ? io_dataIn_0 : _GEN_12; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_45 = 5'h1 == io_wptr_0 ? io_dataIn_0 : _GEN_13; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_46 = 5'h2 == io_wptr_0 ? io_dataIn_0 : _GEN_14; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_47 = 5'h3 == io_wptr_0 ? io_dataIn_0 : _GEN_15; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_48 = 5'h4 == io_wptr_0 ? io_dataIn_0 : _GEN_16; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_49 = 5'h5 == io_wptr_0 ? io_dataIn_0 : _GEN_17; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_50 = 5'h6 == io_wptr_0 ? io_dataIn_0 : _GEN_18; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_51 = 5'h7 == io_wptr_0 ? io_dataIn_0 : _GEN_19; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_52 = 5'h8 == io_wptr_0 ? io_dataIn_0 : _GEN_20; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_53 = 5'h9 == io_wptr_0 ? io_dataIn_0 : _GEN_21; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_54 = 5'ha == io_wptr_0 ? io_dataIn_0 : _GEN_22; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_55 = 5'hb == io_wptr_0 ? io_dataIn_0 : _GEN_23; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_56 = 5'hc == io_wptr_0 ? io_dataIn_0 : _GEN_24; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_57 = 5'hd == io_wptr_0 ? io_dataIn_0 : _GEN_25; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_58 = 5'he == io_wptr_0 ? io_dataIn_0 : _GEN_26; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_59 = 5'hf == io_wptr_0 ? io_dataIn_0 : _GEN_27; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_60 = 5'h10 == io_wptr_0 ? io_dataIn_0 : _GEN_28; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_61 = 5'h11 == io_wptr_0 ? io_dataIn_0 : _GEN_29; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_62 = 5'h12 == io_wptr_0 ? io_dataIn_0 : _GEN_30; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_63 = 5'h13 == io_wptr_0 ? io_dataIn_0 : _GEN_31; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_64 = 5'h14 == io_wptr_0 ? io_dataIn_0 : _GEN_32; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_65 = 5'h15 == io_wptr_0 ? io_dataIn_0 : _GEN_33; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_66 = 5'h16 == io_wptr_0 ? io_dataIn_0 : _GEN_34; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_67 = 5'h17 == io_wptr_0 ? io_dataIn_0 : _GEN_35; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_68 = 5'h18 == io_wptr_0 ? io_dataIn_0 : _GEN_36; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_69 = 5'h19 == io_wptr_0 ? io_dataIn_0 : _GEN_37; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_70 = 5'h1a == io_wptr_0 ? io_dataIn_0 : _GEN_38; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_71 = 5'h1b == io_wptr_0 ? io_dataIn_0 : _GEN_39; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_72 = 5'h1c == io_wptr_0 ? io_dataIn_0 : _GEN_40; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_73 = 5'h1d == io_wptr_0 ? io_dataIn_0 : _GEN_41; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_74 = 5'h1e == io_wptr_0 ? io_dataIn_0 : _GEN_42; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_75 = 5'h1f == io_wptr_0 ? io_dataIn_0 : _GEN_43; // @[util.scala 72:23 util.scala 72:23]
  wire [31:0] _GEN_204 = 5'h0 == io_wptr_1 ? io_dataIn_1 : _GEN_12; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_205 = 5'h1 == io_wptr_1 ? io_dataIn_1 : _GEN_13; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_206 = 5'h2 == io_wptr_1 ? io_dataIn_1 : _GEN_14; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_207 = 5'h3 == io_wptr_1 ? io_dataIn_1 : _GEN_15; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_208 = 5'h4 == io_wptr_1 ? io_dataIn_1 : _GEN_16; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_209 = 5'h5 == io_wptr_1 ? io_dataIn_1 : _GEN_17; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_210 = 5'h6 == io_wptr_1 ? io_dataIn_1 : _GEN_18; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_211 = 5'h7 == io_wptr_1 ? io_dataIn_1 : _GEN_19; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_212 = 5'h8 == io_wptr_1 ? io_dataIn_1 : _GEN_20; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_213 = 5'h9 == io_wptr_1 ? io_dataIn_1 : _GEN_21; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_214 = 5'ha == io_wptr_1 ? io_dataIn_1 : _GEN_22; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_215 = 5'hb == io_wptr_1 ? io_dataIn_1 : _GEN_23; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_216 = 5'hc == io_wptr_1 ? io_dataIn_1 : _GEN_24; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_217 = 5'hd == io_wptr_1 ? io_dataIn_1 : _GEN_25; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_218 = 5'he == io_wptr_1 ? io_dataIn_1 : _GEN_26; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_219 = 5'hf == io_wptr_1 ? io_dataIn_1 : _GEN_27; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_220 = 5'h10 == io_wptr_1 ? io_dataIn_1 : _GEN_28; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_221 = 5'h11 == io_wptr_1 ? io_dataIn_1 : _GEN_29; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_222 = 5'h12 == io_wptr_1 ? io_dataIn_1 : _GEN_30; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_223 = 5'h13 == io_wptr_1 ? io_dataIn_1 : _GEN_31; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_224 = 5'h14 == io_wptr_1 ? io_dataIn_1 : _GEN_32; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_225 = 5'h15 == io_wptr_1 ? io_dataIn_1 : _GEN_33; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_226 = 5'h16 == io_wptr_1 ? io_dataIn_1 : _GEN_34; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_227 = 5'h17 == io_wptr_1 ? io_dataIn_1 : _GEN_35; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_228 = 5'h18 == io_wptr_1 ? io_dataIn_1 : _GEN_36; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_229 = 5'h19 == io_wptr_1 ? io_dataIn_1 : _GEN_37; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_230 = 5'h1a == io_wptr_1 ? io_dataIn_1 : _GEN_38; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_231 = 5'h1b == io_wptr_1 ? io_dataIn_1 : _GEN_39; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_232 = 5'h1c == io_wptr_1 ? io_dataIn_1 : _GEN_40; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_233 = 5'h1d == io_wptr_1 ? io_dataIn_1 : _GEN_41; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_234 = 5'h1e == io_wptr_1 ? io_dataIn_1 : _GEN_42; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_235 = 5'h1f == io_wptr_1 ? io_dataIn_1 : _GEN_43; // @[util.scala 79:23 util.scala 79:23]
  wire [31:0] _GEN_268 = 5'h0 == io_wptr_0 ? io_dataIn_0 : table_0; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_269 = 5'h1 == io_wptr_0 ? io_dataIn_0 : table_1; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_270 = 5'h2 == io_wptr_0 ? io_dataIn_0 : table_2; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_271 = 5'h3 == io_wptr_0 ? io_dataIn_0 : table_3; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_272 = 5'h4 == io_wptr_0 ? io_dataIn_0 : table_4; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_273 = 5'h5 == io_wptr_0 ? io_dataIn_0 : table_5; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_274 = 5'h6 == io_wptr_0 ? io_dataIn_0 : table_6; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_275 = 5'h7 == io_wptr_0 ? io_dataIn_0 : table_7; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_276 = 5'h8 == io_wptr_0 ? io_dataIn_0 : table_8; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_277 = 5'h9 == io_wptr_0 ? io_dataIn_0 : table_9; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_278 = 5'ha == io_wptr_0 ? io_dataIn_0 : table_10; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_279 = 5'hb == io_wptr_0 ? io_dataIn_0 : table_11; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_280 = 5'hc == io_wptr_0 ? io_dataIn_0 : table_12; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_281 = 5'hd == io_wptr_0 ? io_dataIn_0 : table_13; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_282 = 5'he == io_wptr_0 ? io_dataIn_0 : table_14; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_283 = 5'hf == io_wptr_0 ? io_dataIn_0 : table_15; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_284 = 5'h10 == io_wptr_0 ? io_dataIn_0 : table_16; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_285 = 5'h11 == io_wptr_0 ? io_dataIn_0 : table_17; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_286 = 5'h12 == io_wptr_0 ? io_dataIn_0 : table_18; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_287 = 5'h13 == io_wptr_0 ? io_dataIn_0 : table_19; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_288 = 5'h14 == io_wptr_0 ? io_dataIn_0 : table_20; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_289 = 5'h15 == io_wptr_0 ? io_dataIn_0 : table_21; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_290 = 5'h16 == io_wptr_0 ? io_dataIn_0 : table_22; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_291 = 5'h17 == io_wptr_0 ? io_dataIn_0 : table_23; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_292 = 5'h18 == io_wptr_0 ? io_dataIn_0 : table_24; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_293 = 5'h19 == io_wptr_0 ? io_dataIn_0 : table_25; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_294 = 5'h1a == io_wptr_0 ? io_dataIn_0 : table_26; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_295 = 5'h1b == io_wptr_0 ? io_dataIn_0 : table_27; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_296 = 5'h1c == io_wptr_0 ? io_dataIn_0 : table_28; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_297 = 5'h1d == io_wptr_0 ? io_dataIn_0 : table_29; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_298 = 5'h1e == io_wptr_0 ? io_dataIn_0 : table_30; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_299 = 5'h1f == io_wptr_0 ? io_dataIn_0 : table_31; // @[util.scala 83:23 util.scala 83:23 util.scala 16:22]
  wire [31:0] _GEN_300 = 5'h0 == io_wptr_1 ? io_dataIn_1 : _GEN_268; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_301 = 5'h1 == io_wptr_1 ? io_dataIn_1 : _GEN_269; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_302 = 5'h2 == io_wptr_1 ? io_dataIn_1 : _GEN_270; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_303 = 5'h3 == io_wptr_1 ? io_dataIn_1 : _GEN_271; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_304 = 5'h4 == io_wptr_1 ? io_dataIn_1 : _GEN_272; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_305 = 5'h5 == io_wptr_1 ? io_dataIn_1 : _GEN_273; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_306 = 5'h6 == io_wptr_1 ? io_dataIn_1 : _GEN_274; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_307 = 5'h7 == io_wptr_1 ? io_dataIn_1 : _GEN_275; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_308 = 5'h8 == io_wptr_1 ? io_dataIn_1 : _GEN_276; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_309 = 5'h9 == io_wptr_1 ? io_dataIn_1 : _GEN_277; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_310 = 5'ha == io_wptr_1 ? io_dataIn_1 : _GEN_278; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_311 = 5'hb == io_wptr_1 ? io_dataIn_1 : _GEN_279; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_312 = 5'hc == io_wptr_1 ? io_dataIn_1 : _GEN_280; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_313 = 5'hd == io_wptr_1 ? io_dataIn_1 : _GEN_281; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_314 = 5'he == io_wptr_1 ? io_dataIn_1 : _GEN_282; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_315 = 5'hf == io_wptr_1 ? io_dataIn_1 : _GEN_283; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_316 = 5'h10 == io_wptr_1 ? io_dataIn_1 : _GEN_284; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_317 = 5'h11 == io_wptr_1 ? io_dataIn_1 : _GEN_285; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_318 = 5'h12 == io_wptr_1 ? io_dataIn_1 : _GEN_286; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_319 = 5'h13 == io_wptr_1 ? io_dataIn_1 : _GEN_287; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_320 = 5'h14 == io_wptr_1 ? io_dataIn_1 : _GEN_288; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_321 = 5'h15 == io_wptr_1 ? io_dataIn_1 : _GEN_289; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_322 = 5'h16 == io_wptr_1 ? io_dataIn_1 : _GEN_290; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_323 = 5'h17 == io_wptr_1 ? io_dataIn_1 : _GEN_291; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_324 = 5'h18 == io_wptr_1 ? io_dataIn_1 : _GEN_292; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_325 = 5'h19 == io_wptr_1 ? io_dataIn_1 : _GEN_293; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_326 = 5'h1a == io_wptr_1 ? io_dataIn_1 : _GEN_294; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_327 = 5'h1b == io_wptr_1 ? io_dataIn_1 : _GEN_295; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_328 = 5'h1c == io_wptr_1 ? io_dataIn_1 : _GEN_296; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_329 = 5'h1d == io_wptr_1 ? io_dataIn_1 : _GEN_297; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_330 = 5'h1e == io_wptr_1 ? io_dataIn_1 : _GEN_298; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_331 = 5'h1f == io_wptr_1 ? io_dataIn_1 : _GEN_299; // @[util.scala 84:23 util.scala 84:23]
  wire [31:0] _GEN_364 = 5'h0 == io_wptr_1 ? io_dataIn_1 : table_0; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_365 = 5'h1 == io_wptr_1 ? io_dataIn_1 : table_1; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_366 = 5'h2 == io_wptr_1 ? io_dataIn_1 : table_2; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_367 = 5'h3 == io_wptr_1 ? io_dataIn_1 : table_3; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_368 = 5'h4 == io_wptr_1 ? io_dataIn_1 : table_4; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_369 = 5'h5 == io_wptr_1 ? io_dataIn_1 : table_5; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_370 = 5'h6 == io_wptr_1 ? io_dataIn_1 : table_6; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_371 = 5'h7 == io_wptr_1 ? io_dataIn_1 : table_7; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_372 = 5'h8 == io_wptr_1 ? io_dataIn_1 : table_8; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_373 = 5'h9 == io_wptr_1 ? io_dataIn_1 : table_9; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_374 = 5'ha == io_wptr_1 ? io_dataIn_1 : table_10; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_375 = 5'hb == io_wptr_1 ? io_dataIn_1 : table_11; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_376 = 5'hc == io_wptr_1 ? io_dataIn_1 : table_12; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_377 = 5'hd == io_wptr_1 ? io_dataIn_1 : table_13; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_378 = 5'he == io_wptr_1 ? io_dataIn_1 : table_14; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_379 = 5'hf == io_wptr_1 ? io_dataIn_1 : table_15; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_380 = 5'h10 == io_wptr_1 ? io_dataIn_1 : table_16; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_381 = 5'h11 == io_wptr_1 ? io_dataIn_1 : table_17; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_382 = 5'h12 == io_wptr_1 ? io_dataIn_1 : table_18; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_383 = 5'h13 == io_wptr_1 ? io_dataIn_1 : table_19; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_384 = 5'h14 == io_wptr_1 ? io_dataIn_1 : table_20; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_385 = 5'h15 == io_wptr_1 ? io_dataIn_1 : table_21; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_386 = 5'h16 == io_wptr_1 ? io_dataIn_1 : table_22; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_387 = 5'h17 == io_wptr_1 ? io_dataIn_1 : table_23; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_388 = 5'h18 == io_wptr_1 ? io_dataIn_1 : table_24; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_389 = 5'h19 == io_wptr_1 ? io_dataIn_1 : table_25; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_390 = 5'h1a == io_wptr_1 ? io_dataIn_1 : table_26; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_391 = 5'h1b == io_wptr_1 ? io_dataIn_1 : table_27; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_392 = 5'h1c == io_wptr_1 ? io_dataIn_1 : table_28; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_393 = 5'h1d == io_wptr_1 ? io_dataIn_1 : table_29; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_394 = 5'h1e == io_wptr_1 ? io_dataIn_1 : table_30; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_395 = 5'h1f == io_wptr_1 ? io_dataIn_1 : table_31; // @[util.scala 88:23 util.scala 88:23 util.scala 16:22]
  wire [31:0] _GEN_396 = io_writeFlag_1 ? _GEN_364 : table_0; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_397 = io_writeFlag_1 ? _GEN_365 : table_1; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_398 = io_writeFlag_1 ? _GEN_366 : table_2; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_399 = io_writeFlag_1 ? _GEN_367 : table_3; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_400 = io_writeFlag_1 ? _GEN_368 : table_4; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_401 = io_writeFlag_1 ? _GEN_369 : table_5; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_402 = io_writeFlag_1 ? _GEN_370 : table_6; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_403 = io_writeFlag_1 ? _GEN_371 : table_7; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_404 = io_writeFlag_1 ? _GEN_372 : table_8; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_405 = io_writeFlag_1 ? _GEN_373 : table_9; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_406 = io_writeFlag_1 ? _GEN_374 : table_10; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_407 = io_writeFlag_1 ? _GEN_375 : table_11; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_408 = io_writeFlag_1 ? _GEN_376 : table_12; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_409 = io_writeFlag_1 ? _GEN_377 : table_13; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_410 = io_writeFlag_1 ? _GEN_378 : table_14; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_411 = io_writeFlag_1 ? _GEN_379 : table_15; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_412 = io_writeFlag_1 ? _GEN_380 : table_16; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_413 = io_writeFlag_1 ? _GEN_381 : table_17; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_414 = io_writeFlag_1 ? _GEN_382 : table_18; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_415 = io_writeFlag_1 ? _GEN_383 : table_19; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_416 = io_writeFlag_1 ? _GEN_384 : table_20; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_417 = io_writeFlag_1 ? _GEN_385 : table_21; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_418 = io_writeFlag_1 ? _GEN_386 : table_22; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_419 = io_writeFlag_1 ? _GEN_387 : table_23; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_420 = io_writeFlag_1 ? _GEN_388 : table_24; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_421 = io_writeFlag_1 ? _GEN_389 : table_25; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_422 = io_writeFlag_1 ? _GEN_390 : table_26; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_423 = io_writeFlag_1 ? _GEN_391 : table_27; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_424 = io_writeFlag_1 ? _GEN_392 : table_28; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_425 = io_writeFlag_1 ? _GEN_393 : table_29; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_426 = io_writeFlag_1 ? _GEN_394 : table_30; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_427 = io_writeFlag_1 ? _GEN_395 : table_31; // @[util.scala 87:30 util.scala 16:22]
  wire [31:0] _GEN_428 = io_writeFlag_0 ? _GEN_268 : _GEN_396; // @[util.scala 85:30]
  wire [31:0] _GEN_429 = io_writeFlag_0 ? _GEN_269 : _GEN_397; // @[util.scala 85:30]
  wire [31:0] _GEN_430 = io_writeFlag_0 ? _GEN_270 : _GEN_398; // @[util.scala 85:30]
  wire [31:0] _GEN_431 = io_writeFlag_0 ? _GEN_271 : _GEN_399; // @[util.scala 85:30]
  wire [31:0] _GEN_432 = io_writeFlag_0 ? _GEN_272 : _GEN_400; // @[util.scala 85:30]
  wire [31:0] _GEN_433 = io_writeFlag_0 ? _GEN_273 : _GEN_401; // @[util.scala 85:30]
  wire [31:0] _GEN_434 = io_writeFlag_0 ? _GEN_274 : _GEN_402; // @[util.scala 85:30]
  wire [31:0] _GEN_435 = io_writeFlag_0 ? _GEN_275 : _GEN_403; // @[util.scala 85:30]
  wire [31:0] _GEN_436 = io_writeFlag_0 ? _GEN_276 : _GEN_404; // @[util.scala 85:30]
  wire [31:0] _GEN_437 = io_writeFlag_0 ? _GEN_277 : _GEN_405; // @[util.scala 85:30]
  wire [31:0] _GEN_438 = io_writeFlag_0 ? _GEN_278 : _GEN_406; // @[util.scala 85:30]
  wire [31:0] _GEN_439 = io_writeFlag_0 ? _GEN_279 : _GEN_407; // @[util.scala 85:30]
  wire [31:0] _GEN_440 = io_writeFlag_0 ? _GEN_280 : _GEN_408; // @[util.scala 85:30]
  wire [31:0] _GEN_441 = io_writeFlag_0 ? _GEN_281 : _GEN_409; // @[util.scala 85:30]
  wire [31:0] _GEN_442 = io_writeFlag_0 ? _GEN_282 : _GEN_410; // @[util.scala 85:30]
  wire [31:0] _GEN_443 = io_writeFlag_0 ? _GEN_283 : _GEN_411; // @[util.scala 85:30]
  wire [31:0] _GEN_444 = io_writeFlag_0 ? _GEN_284 : _GEN_412; // @[util.scala 85:30]
  wire [31:0] _GEN_445 = io_writeFlag_0 ? _GEN_285 : _GEN_413; // @[util.scala 85:30]
  wire [31:0] _GEN_446 = io_writeFlag_0 ? _GEN_286 : _GEN_414; // @[util.scala 85:30]
  wire [31:0] _GEN_447 = io_writeFlag_0 ? _GEN_287 : _GEN_415; // @[util.scala 85:30]
  wire [31:0] _GEN_448 = io_writeFlag_0 ? _GEN_288 : _GEN_416; // @[util.scala 85:30]
  wire [31:0] _GEN_449 = io_writeFlag_0 ? _GEN_289 : _GEN_417; // @[util.scala 85:30]
  wire [31:0] _GEN_450 = io_writeFlag_0 ? _GEN_290 : _GEN_418; // @[util.scala 85:30]
  wire [31:0] _GEN_451 = io_writeFlag_0 ? _GEN_291 : _GEN_419; // @[util.scala 85:30]
  wire [31:0] _GEN_452 = io_writeFlag_0 ? _GEN_292 : _GEN_420; // @[util.scala 85:30]
  wire [31:0] _GEN_453 = io_writeFlag_0 ? _GEN_293 : _GEN_421; // @[util.scala 85:30]
  wire [31:0] _GEN_454 = io_writeFlag_0 ? _GEN_294 : _GEN_422; // @[util.scala 85:30]
  wire [31:0] _GEN_455 = io_writeFlag_0 ? _GEN_295 : _GEN_423; // @[util.scala 85:30]
  wire [31:0] _GEN_456 = io_writeFlag_0 ? _GEN_296 : _GEN_424; // @[util.scala 85:30]
  wire [31:0] _GEN_457 = io_writeFlag_0 ? _GEN_297 : _GEN_425; // @[util.scala 85:30]
  wire [31:0] _GEN_458 = io_writeFlag_0 ? _GEN_298 : _GEN_426; // @[util.scala 85:30]
  wire [31:0] _GEN_459 = io_writeFlag_0 ? _GEN_299 : _GEN_427; // @[util.scala 85:30]
  wire [31:0] _GEN_460 = _T_7 ? _GEN_300 : _GEN_428; // @[util.scala 82:39]
  wire [31:0] _GEN_461 = _T_7 ? _GEN_301 : _GEN_429; // @[util.scala 82:39]
  wire [31:0] _GEN_462 = _T_7 ? _GEN_302 : _GEN_430; // @[util.scala 82:39]
  wire [31:0] _GEN_463 = _T_7 ? _GEN_303 : _GEN_431; // @[util.scala 82:39]
  wire [31:0] _GEN_464 = _T_7 ? _GEN_304 : _GEN_432; // @[util.scala 82:39]
  wire [31:0] _GEN_465 = _T_7 ? _GEN_305 : _GEN_433; // @[util.scala 82:39]
  wire [31:0] _GEN_466 = _T_7 ? _GEN_306 : _GEN_434; // @[util.scala 82:39]
  wire [31:0] _GEN_467 = _T_7 ? _GEN_307 : _GEN_435; // @[util.scala 82:39]
  wire [31:0] _GEN_468 = _T_7 ? _GEN_308 : _GEN_436; // @[util.scala 82:39]
  wire [31:0] _GEN_469 = _T_7 ? _GEN_309 : _GEN_437; // @[util.scala 82:39]
  wire [31:0] _GEN_470 = _T_7 ? _GEN_310 : _GEN_438; // @[util.scala 82:39]
  wire [31:0] _GEN_471 = _T_7 ? _GEN_311 : _GEN_439; // @[util.scala 82:39]
  wire [31:0] _GEN_472 = _T_7 ? _GEN_312 : _GEN_440; // @[util.scala 82:39]
  wire [31:0] _GEN_473 = _T_7 ? _GEN_313 : _GEN_441; // @[util.scala 82:39]
  wire [31:0] _GEN_474 = _T_7 ? _GEN_314 : _GEN_442; // @[util.scala 82:39]
  wire [31:0] _GEN_475 = _T_7 ? _GEN_315 : _GEN_443; // @[util.scala 82:39]
  wire [31:0] _GEN_476 = _T_7 ? _GEN_316 : _GEN_444; // @[util.scala 82:39]
  wire [31:0] _GEN_477 = _T_7 ? _GEN_317 : _GEN_445; // @[util.scala 82:39]
  wire [31:0] _GEN_478 = _T_7 ? _GEN_318 : _GEN_446; // @[util.scala 82:39]
  wire [31:0] _GEN_479 = _T_7 ? _GEN_319 : _GEN_447; // @[util.scala 82:39]
  wire [31:0] _GEN_480 = _T_7 ? _GEN_320 : _GEN_448; // @[util.scala 82:39]
  wire [31:0] _GEN_481 = _T_7 ? _GEN_321 : _GEN_449; // @[util.scala 82:39]
  wire [31:0] _GEN_482 = _T_7 ? _GEN_322 : _GEN_450; // @[util.scala 82:39]
  wire [31:0] _GEN_483 = _T_7 ? _GEN_323 : _GEN_451; // @[util.scala 82:39]
  wire [31:0] _GEN_484 = _T_7 ? _GEN_324 : _GEN_452; // @[util.scala 82:39]
  wire [31:0] _GEN_485 = _T_7 ? _GEN_325 : _GEN_453; // @[util.scala 82:39]
  wire [31:0] _GEN_486 = _T_7 ? _GEN_326 : _GEN_454; // @[util.scala 82:39]
  wire [31:0] _GEN_487 = _T_7 ? _GEN_327 : _GEN_455; // @[util.scala 82:39]
  wire [31:0] _GEN_488 = _T_7 ? _GEN_328 : _GEN_456; // @[util.scala 82:39]
  wire [31:0] _GEN_489 = _T_7 ? _GEN_329 : _GEN_457; // @[util.scala 82:39]
  wire [31:0] _GEN_490 = _T_7 ? _GEN_330 : _GEN_458; // @[util.scala 82:39]
  wire [31:0] _GEN_491 = _T_7 ? _GEN_331 : _GEN_459; // @[util.scala 82:39]
  wire [31:0] _GEN_492 = wvalid ? _GEN_12 : _GEN_460; // @[util.scala 80:21]
  wire [31:0] _GEN_493 = wvalid ? _GEN_13 : _GEN_461; // @[util.scala 80:21]
  wire [31:0] _GEN_494 = wvalid ? _GEN_14 : _GEN_462; // @[util.scala 80:21]
  wire [31:0] _GEN_495 = wvalid ? _GEN_15 : _GEN_463; // @[util.scala 80:21]
  wire [31:0] _GEN_496 = wvalid ? _GEN_16 : _GEN_464; // @[util.scala 80:21]
  wire [31:0] _GEN_497 = wvalid ? _GEN_17 : _GEN_465; // @[util.scala 80:21]
  wire [31:0] _GEN_498 = wvalid ? _GEN_18 : _GEN_466; // @[util.scala 80:21]
  wire [31:0] _GEN_499 = wvalid ? _GEN_19 : _GEN_467; // @[util.scala 80:21]
  wire [31:0] _GEN_500 = wvalid ? _GEN_20 : _GEN_468; // @[util.scala 80:21]
  wire [31:0] _GEN_501 = wvalid ? _GEN_21 : _GEN_469; // @[util.scala 80:21]
  wire [31:0] _GEN_502 = wvalid ? _GEN_22 : _GEN_470; // @[util.scala 80:21]
  wire [31:0] _GEN_503 = wvalid ? _GEN_23 : _GEN_471; // @[util.scala 80:21]
  wire [31:0] _GEN_504 = wvalid ? _GEN_24 : _GEN_472; // @[util.scala 80:21]
  wire [31:0] _GEN_505 = wvalid ? _GEN_25 : _GEN_473; // @[util.scala 80:21]
  wire [31:0] _GEN_506 = wvalid ? _GEN_26 : _GEN_474; // @[util.scala 80:21]
  wire [31:0] _GEN_507 = wvalid ? _GEN_27 : _GEN_475; // @[util.scala 80:21]
  wire [31:0] _GEN_508 = wvalid ? _GEN_28 : _GEN_476; // @[util.scala 80:21]
  wire [31:0] _GEN_509 = wvalid ? _GEN_29 : _GEN_477; // @[util.scala 80:21]
  wire [31:0] _GEN_510 = wvalid ? _GEN_30 : _GEN_478; // @[util.scala 80:21]
  wire [31:0] _GEN_511 = wvalid ? _GEN_31 : _GEN_479; // @[util.scala 80:21]
  wire [31:0] _GEN_512 = wvalid ? _GEN_32 : _GEN_480; // @[util.scala 80:21]
  wire [31:0] _GEN_513 = wvalid ? _GEN_33 : _GEN_481; // @[util.scala 80:21]
  wire [31:0] _GEN_514 = wvalid ? _GEN_34 : _GEN_482; // @[util.scala 80:21]
  wire [31:0] _GEN_515 = wvalid ? _GEN_35 : _GEN_483; // @[util.scala 80:21]
  wire [31:0] _GEN_516 = wvalid ? _GEN_36 : _GEN_484; // @[util.scala 80:21]
  wire [31:0] _GEN_517 = wvalid ? _GEN_37 : _GEN_485; // @[util.scala 80:21]
  wire [31:0] _GEN_518 = wvalid ? _GEN_38 : _GEN_486; // @[util.scala 80:21]
  wire [31:0] _GEN_519 = wvalid ? _GEN_39 : _GEN_487; // @[util.scala 80:21]
  wire [31:0] _GEN_520 = wvalid ? _GEN_40 : _GEN_488; // @[util.scala 80:21]
  wire [31:0] _GEN_521 = wvalid ? _GEN_41 : _GEN_489; // @[util.scala 80:21]
  wire [31:0] _GEN_522 = wvalid ? _GEN_42 : _GEN_490; // @[util.scala 80:21]
  wire [31:0] _GEN_523 = wvalid ? _GEN_43 : _GEN_491; // @[util.scala 80:21]
  reg [4:0] eraddr; // @[util.scala 92:19]
  wire [31:0] _GEN_622 = 5'h1 == eraddr ? table_1 : table_0; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_623 = 5'h2 == eraddr ? table_2 : _GEN_622; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_624 = 5'h3 == eraddr ? table_3 : _GEN_623; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_625 = 5'h4 == eraddr ? table_4 : _GEN_624; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_626 = 5'h5 == eraddr ? table_5 : _GEN_625; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_627 = 5'h6 == eraddr ? table_6 : _GEN_626; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_628 = 5'h7 == eraddr ? table_7 : _GEN_627; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_629 = 5'h8 == eraddr ? table_8 : _GEN_628; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_630 = 5'h9 == eraddr ? table_9 : _GEN_629; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_631 = 5'ha == eraddr ? table_10 : _GEN_630; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_632 = 5'hb == eraddr ? table_11 : _GEN_631; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_633 = 5'hc == eraddr ? table_12 : _GEN_632; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_634 = 5'hd == eraddr ? table_13 : _GEN_633; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_635 = 5'he == eraddr ? table_14 : _GEN_634; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_636 = 5'hf == eraddr ? table_15 : _GEN_635; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_637 = 5'h10 == eraddr ? table_16 : _GEN_636; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_638 = 5'h11 == eraddr ? table_17 : _GEN_637; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_639 = 5'h12 == eraddr ? table_18 : _GEN_638; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_640 = 5'h13 == eraddr ? table_19 : _GEN_639; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_641 = 5'h14 == eraddr ? table_20 : _GEN_640; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_642 = 5'h15 == eraddr ? table_21 : _GEN_641; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_643 = 5'h16 == eraddr ? table_22 : _GEN_642; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_644 = 5'h17 == eraddr ? table_23 : _GEN_643; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_645 = 5'h18 == eraddr ? table_24 : _GEN_644; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_646 = 5'h19 == eraddr ? table_25 : _GEN_645; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_647 = 5'h1a == eraddr ? table_26 : _GEN_646; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_648 = 5'h1b == eraddr ? table_27 : _GEN_647; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_649 = 5'h1c == eraddr ? table_28 : _GEN_648; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_650 = 5'h1d == eraddr ? table_29 : _GEN_649; // @[util.scala 99:16 util.scala 99:16]
  wire [31:0] _GEN_651 = 5'h1e == eraddr ? table_30 : _GEN_650; // @[util.scala 99:16 util.scala 99:16]
  assign io_data_0 = table_0; // @[util.scala 53:11]
  assign io_data_1 = table_1; // @[util.scala 53:11]
  assign io_data_2 = table_2; // @[util.scala 53:11]
  assign io_data_3 = table_3; // @[util.scala 53:11]
  assign io_data_4 = table_4; // @[util.scala 53:11]
  assign io_data_5 = table_5; // @[util.scala 53:11]
  assign io_data_6 = table_6; // @[util.scala 53:11]
  assign io_data_7 = table_7; // @[util.scala 53:11]
  assign io_data_8 = table_8; // @[util.scala 53:11]
  assign io_data_9 = table_9; // @[util.scala 53:11]
  assign io_data_10 = table_10; // @[util.scala 53:11]
  assign io_data_11 = table_11; // @[util.scala 53:11]
  assign io_data_12 = table_12; // @[util.scala 53:11]
  assign io_data_13 = table_13; // @[util.scala 53:11]
  assign io_data_16 = table_16; // @[util.scala 53:11]
  assign io_data_17 = table_17; // @[util.scala 53:11]
  assign io_data_18 = table_18; // @[util.scala 53:11]
  assign config_awready = status == 3'h0; // @[util.scala 55:28]
  assign config_arready = status == 3'h0; // @[util.scala 56:28]
  assign config_wready = status == 3'h1; // @[util.scala 54:27]
  assign config_rdata = 5'h1f == eraddr ? table_31 : _GEN_651; // @[util.scala 99:16 util.scala 99:16]
  assign config_rvalid = status == 3'h5; // @[util.scala 57:27]
  assign config_bvalid = status == 3'h3; // @[util.scala 58:27]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 16:22]
      table_0 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h0 == io_wptr_1) begin // @[util.scala 73:23]
        table_0 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_0 <= _GEN_44;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_0 <= _GEN_44;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_0 <= _GEN_204;
    end else begin
      table_0 <= _GEN_492;
    end
    if (reset) begin // @[util.scala 16:22]
      table_1 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1 == io_wptr_1) begin // @[util.scala 73:23]
        table_1 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_1 <= _GEN_45;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_1 <= _GEN_45;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_1 <= _GEN_205;
    end else begin
      table_1 <= _GEN_493;
    end
    if (reset) begin // @[util.scala 16:22]
      table_2 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h2 == io_wptr_1) begin // @[util.scala 73:23]
        table_2 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_2 <= _GEN_46;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_2 <= _GEN_46;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_2 <= _GEN_206;
    end else begin
      table_2 <= _GEN_494;
    end
    if (reset) begin // @[util.scala 16:22]
      table_3 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h3 == io_wptr_1) begin // @[util.scala 73:23]
        table_3 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_3 <= _GEN_47;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_3 <= _GEN_47;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_3 <= _GEN_207;
    end else begin
      table_3 <= _GEN_495;
    end
    if (reset) begin // @[util.scala 16:22]
      table_4 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h4 == io_wptr_1) begin // @[util.scala 73:23]
        table_4 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_4 <= _GEN_48;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_4 <= _GEN_48;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_4 <= _GEN_208;
    end else begin
      table_4 <= _GEN_496;
    end
    if (reset) begin // @[util.scala 16:22]
      table_5 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h5 == io_wptr_1) begin // @[util.scala 73:23]
        table_5 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_5 <= _GEN_49;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_5 <= _GEN_49;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_5 <= _GEN_209;
    end else begin
      table_5 <= _GEN_497;
    end
    if (reset) begin // @[util.scala 16:22]
      table_6 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h6 == io_wptr_1) begin // @[util.scala 73:23]
        table_6 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_6 <= _GEN_50;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_6 <= _GEN_50;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_6 <= _GEN_210;
    end else begin
      table_6 <= _GEN_498;
    end
    if (reset) begin // @[util.scala 16:22]
      table_7 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h7 == io_wptr_1) begin // @[util.scala 73:23]
        table_7 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_7 <= _GEN_51;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_7 <= _GEN_51;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_7 <= _GEN_211;
    end else begin
      table_7 <= _GEN_499;
    end
    if (reset) begin // @[util.scala 16:22]
      table_8 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h8 == io_wptr_1) begin // @[util.scala 73:23]
        table_8 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_8 <= _GEN_52;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_8 <= _GEN_52;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_8 <= _GEN_212;
    end else begin
      table_8 <= _GEN_500;
    end
    if (reset) begin // @[util.scala 16:22]
      table_9 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h9 == io_wptr_1) begin // @[util.scala 73:23]
        table_9 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_9 <= _GEN_53;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_9 <= _GEN_53;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_9 <= _GEN_213;
    end else begin
      table_9 <= _GEN_501;
    end
    if (reset) begin // @[util.scala 16:22]
      table_10 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'ha == io_wptr_1) begin // @[util.scala 73:23]
        table_10 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_10 <= _GEN_54;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_10 <= _GEN_54;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_10 <= _GEN_214;
    end else begin
      table_10 <= _GEN_502;
    end
    if (reset) begin // @[util.scala 16:22]
      table_11 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hb == io_wptr_1) begin // @[util.scala 73:23]
        table_11 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_11 <= _GEN_55;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_11 <= _GEN_55;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_11 <= _GEN_215;
    end else begin
      table_11 <= _GEN_503;
    end
    if (reset) begin // @[util.scala 16:22]
      table_12 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hc == io_wptr_1) begin // @[util.scala 73:23]
        table_12 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_12 <= _GEN_56;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_12 <= _GEN_56;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_12 <= _GEN_216;
    end else begin
      table_12 <= _GEN_504;
    end
    if (reset) begin // @[util.scala 16:22]
      table_13 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hd == io_wptr_1) begin // @[util.scala 73:23]
        table_13 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_13 <= _GEN_57;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_13 <= _GEN_57;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_13 <= _GEN_217;
    end else begin
      table_13 <= _GEN_505;
    end
    if (reset) begin // @[util.scala 16:22]
      table_14 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'he == io_wptr_1) begin // @[util.scala 73:23]
        table_14 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_14 <= _GEN_58;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_14 <= _GEN_58;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_14 <= _GEN_218;
    end else begin
      table_14 <= _GEN_506;
    end
    if (reset) begin // @[util.scala 16:22]
      table_15 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'hf == io_wptr_1) begin // @[util.scala 73:23]
        table_15 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_15 <= _GEN_59;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_15 <= _GEN_59;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_15 <= _GEN_219;
    end else begin
      table_15 <= _GEN_507;
    end
    if (reset) begin // @[util.scala 16:22]
      table_16 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h10 == io_wptr_1) begin // @[util.scala 73:23]
        table_16 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_16 <= _GEN_60;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_16 <= _GEN_60;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_16 <= _GEN_220;
    end else begin
      table_16 <= _GEN_508;
    end
    if (reset) begin // @[util.scala 16:22]
      table_17 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h11 == io_wptr_1) begin // @[util.scala 73:23]
        table_17 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_17 <= _GEN_61;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_17 <= _GEN_61;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_17 <= _GEN_221;
    end else begin
      table_17 <= _GEN_509;
    end
    if (reset) begin // @[util.scala 16:22]
      table_18 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h12 == io_wptr_1) begin // @[util.scala 73:23]
        table_18 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_18 <= _GEN_62;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_18 <= _GEN_62;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_18 <= _GEN_222;
    end else begin
      table_18 <= _GEN_510;
    end
    if (reset) begin // @[util.scala 16:22]
      table_19 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h13 == io_wptr_1) begin // @[util.scala 73:23]
        table_19 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_19 <= _GEN_63;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_19 <= _GEN_63;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_19 <= _GEN_223;
    end else begin
      table_19 <= _GEN_511;
    end
    if (reset) begin // @[util.scala 16:22]
      table_20 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h14 == io_wptr_1) begin // @[util.scala 73:23]
        table_20 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_20 <= _GEN_64;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_20 <= _GEN_64;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_20 <= _GEN_224;
    end else begin
      table_20 <= _GEN_512;
    end
    if (reset) begin // @[util.scala 16:22]
      table_21 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h15 == io_wptr_1) begin // @[util.scala 73:23]
        table_21 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_21 <= _GEN_65;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_21 <= _GEN_65;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_21 <= _GEN_225;
    end else begin
      table_21 <= _GEN_513;
    end
    if (reset) begin // @[util.scala 16:22]
      table_22 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h16 == io_wptr_1) begin // @[util.scala 73:23]
        table_22 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_22 <= _GEN_66;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_22 <= _GEN_66;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_22 <= _GEN_226;
    end else begin
      table_22 <= _GEN_514;
    end
    if (reset) begin // @[util.scala 16:22]
      table_23 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h17 == io_wptr_1) begin // @[util.scala 73:23]
        table_23 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_23 <= _GEN_67;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_23 <= _GEN_67;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_23 <= _GEN_227;
    end else begin
      table_23 <= _GEN_515;
    end
    if (reset) begin // @[util.scala 16:22]
      table_24 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h18 == io_wptr_1) begin // @[util.scala 73:23]
        table_24 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_24 <= _GEN_68;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_24 <= _GEN_68;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_24 <= _GEN_228;
    end else begin
      table_24 <= _GEN_516;
    end
    if (reset) begin // @[util.scala 16:22]
      table_25 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h19 == io_wptr_1) begin // @[util.scala 73:23]
        table_25 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_25 <= _GEN_69;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_25 <= _GEN_69;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_25 <= _GEN_229;
    end else begin
      table_25 <= _GEN_517;
    end
    if (reset) begin // @[util.scala 16:22]
      table_26 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1a == io_wptr_1) begin // @[util.scala 73:23]
        table_26 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_26 <= _GEN_70;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_26 <= _GEN_70;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_26 <= _GEN_230;
    end else begin
      table_26 <= _GEN_518;
    end
    if (reset) begin // @[util.scala 16:22]
      table_27 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1b == io_wptr_1) begin // @[util.scala 73:23]
        table_27 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_27 <= _GEN_71;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_27 <= _GEN_71;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_27 <= _GEN_231;
    end else begin
      table_27 <= _GEN_519;
    end
    if (reset) begin // @[util.scala 16:22]
      table_28 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1c == io_wptr_1) begin // @[util.scala 73:23]
        table_28 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_28 <= _GEN_72;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_28 <= _GEN_72;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_28 <= _GEN_232;
    end else begin
      table_28 <= _GEN_520;
    end
    if (reset) begin // @[util.scala 16:22]
      table_29 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1d == io_wptr_1) begin // @[util.scala 73:23]
        table_29 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_29 <= _GEN_73;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_29 <= _GEN_73;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_29 <= _GEN_233;
    end else begin
      table_29 <= _GEN_521;
    end
    if (reset) begin // @[util.scala 16:22]
      table_30 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1e == io_wptr_1) begin // @[util.scala 73:23]
        table_30 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_30 <= _GEN_74;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_30 <= _GEN_74;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_30 <= _GEN_234;
    end else begin
      table_30 <= _GEN_522;
    end
    if (reset) begin // @[util.scala 16:22]
      table_31 <= 32'h0; // @[util.scala 16:22]
    end else if (wvalid & (io_writeFlag_0 & io_writeFlag_1)) begin // @[util.scala 70:43]
      if (5'h1f == io_wptr_1) begin // @[util.scala 73:23]
        table_31 <= io_dataIn_1; // @[util.scala 73:23]
      end else begin
        table_31 <= _GEN_75;
      end
    end else if (wvalid & io_writeFlag_0) begin // @[util.scala 74:40]
      table_31 <= _GEN_75;
    end else if (wvalid & io_writeFlag_1) begin // @[util.scala 77:40]
      table_31 <= _GEN_235;
    end else begin
      table_31 <= _GEN_523;
    end
    if (reset) begin // @[util.scala 26:23]
      status <= 3'h0; // @[util.scala 26:23]
    end else if (status == 3'h0) begin // @[util.scala 28:28]
      if (config_awvalid) begin // @[util.scala 29:25]
        status <= 3'h1; // @[util.scala 30:14]
      end else if (config_arvalid) begin // @[util.scala 31:31]
        status <= 3'h4; // @[util.scala 32:14]
      end
    end else if (status == 3'h1) begin // @[util.scala 34:35]
      if (config_wvalid) begin // @[util.scala 35:24]
        status <= 3'h2; // @[util.scala 36:14]
      end
    end else if (status == 3'h2) begin // @[util.scala 38:34]
      status <= 3'h3; // @[util.scala 39:12]
    end else begin
      status <= _GEN_7;
    end
    if (config_awvalid & config_awready) begin // @[util.scala 66:41]
      ewaddr <= config_awaddr[6:2]; // @[util.scala 67:12]
    end
    if (config_arvalid & config_arready) begin // @[util.scala 93:41]
      eraddr <= config_araddr[6:2]; // @[util.scala 94:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  table_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  table_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  table_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  table_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  table_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  table_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  table_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  table_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  table_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  table_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  table_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  table_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  table_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  table_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  table_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  table_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  table_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  table_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  table_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  table_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  table_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  table_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  table_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  table_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  table_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  table_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  table_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  table_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  table_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  table_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  table_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  table_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  status = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  ewaddr = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  eraddr = _RAND_34[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module controller(
  input         clock,
  input         reset,
  output [31:0] io_data_0,
  output [31:0] io_data_1,
  output [31:0] io_data_2,
  output [31:0] io_data_3,
  output [31:0] io_data_4,
  output [31:0] io_data_5,
  output [31:0] io_data_6,
  output [31:0] io_data_7,
  output [31:0] io_data_8,
  output [31:0] io_data_9,
  output [31:0] io_data_10,
  output [31:0] io_data_11,
  output [31:0] io_data_16,
  output [31:0] io_data_17,
  output [31:0] io_data_18,
  input         io_fin_0,
  input         io_fin_1,
  input         io_fin_2,
  input         io_fin_3,
  input         io_fin_4,
  input         io_fin_5,
  input         io_fin_6,
  input         io_fin_7,
  input         io_fin_8,
  input         io_fin_9,
  input         io_fin_10,
  input         io_fin_11,
  input         io_fin_12,
  input         io_fin_13,
  input         io_fin_14,
  input         io_fin_15,
  input         io_fin_16,
  output        io_signal,
  output        io_start,
  output [31:0] io_level,
  input  [31:0] io_unvisited_size,
  input  [63:0] io_traveled_edges,
  input  [63:0] io_config_awaddr,
  input         io_config_awvalid,
  output        io_config_awready,
  input  [63:0] io_config_araddr,
  input         io_config_arvalid,
  output        io_config_arready,
  input  [31:0] io_config_wdata,
  input         io_config_wvalid,
  output        io_config_wready,
  output [31:0] io_config_rdata,
  output        io_config_rvalid,
  input         io_config_rready,
  output        io_config_bvalid,
  input         io_config_bready,
  output        io_flush_cache,
  input         io_flush_cache_end,
  input         io_signal_ack,
  input         io_performance_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  controls_clock; // @[BFS.scala 1105:24]
  wire  controls_reset; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_0; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_1; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_2; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_3; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_4; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_5; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_6; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_7; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_8; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_9; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_10; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_11; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_12; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_13; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_16; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_17; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_data_18; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_dataIn_0; // @[BFS.scala 1105:24]
  wire [31:0] controls_io_dataIn_1; // @[BFS.scala 1105:24]
  wire  controls_io_writeFlag_0; // @[BFS.scala 1105:24]
  wire  controls_io_writeFlag_1; // @[BFS.scala 1105:24]
  wire [4:0] controls_io_wptr_0; // @[BFS.scala 1105:24]
  wire [4:0] controls_io_wptr_1; // @[BFS.scala 1105:24]
  wire [63:0] controls_config_awaddr; // @[BFS.scala 1105:24]
  wire  controls_config_awvalid; // @[BFS.scala 1105:24]
  wire  controls_config_awready; // @[BFS.scala 1105:24]
  wire [63:0] controls_config_araddr; // @[BFS.scala 1105:24]
  wire  controls_config_arvalid; // @[BFS.scala 1105:24]
  wire  controls_config_arready; // @[BFS.scala 1105:24]
  wire [31:0] controls_config_wdata; // @[BFS.scala 1105:24]
  wire  controls_config_wvalid; // @[BFS.scala 1105:24]
  wire  controls_config_wready; // @[BFS.scala 1105:24]
  wire [31:0] controls_config_rdata; // @[BFS.scala 1105:24]
  wire  controls_config_rvalid; // @[BFS.scala 1105:24]
  wire  controls_config_rready; // @[BFS.scala 1105:24]
  wire  controls_config_bvalid; // @[BFS.scala 1105:24]
  wire  controls_config_bready; // @[BFS.scala 1105:24]
  (*dont_touch = "true" *)reg [31:0] level; // @[BFS.scala 1106:22]
  (*dont_touch = "true" *)reg [2:0] status; // @[BFS.scala 1116:23]
  wire  start = controls_io_data_0[0] & ~controls_io_data_0[1]; // @[BFS.scala 1117:38]
  reg  FIN_0; // @[BFS.scala 1118:20]
  reg  FIN_1; // @[BFS.scala 1118:20]
  reg  FIN_2; // @[BFS.scala 1118:20]
  reg  FIN_3; // @[BFS.scala 1118:20]
  reg  FIN_4; // @[BFS.scala 1118:20]
  reg  FIN_5; // @[BFS.scala 1118:20]
  reg  FIN_6; // @[BFS.scala 1118:20]
  reg  FIN_7; // @[BFS.scala 1118:20]
  reg  FIN_8; // @[BFS.scala 1118:20]
  reg  FIN_9; // @[BFS.scala 1118:20]
  reg  FIN_10; // @[BFS.scala 1118:20]
  reg  FIN_11; // @[BFS.scala 1118:20]
  reg  FIN_12; // @[BFS.scala 1118:20]
  reg  FIN_13; // @[BFS.scala 1118:20]
  reg  FIN_14; // @[BFS.scala 1118:20]
  reg  FIN_15; // @[BFS.scala 1118:20]
  reg  FIN_16; // @[BFS.scala 1118:20]
  wire [63:0] _new_tep_T = {controls_io_data_12,controls_io_data_13}; // @[Cat.scala 30:58]
  wire [63:0] new_tep = _new_tep_T + io_traveled_edges; // @[BFS.scala 1119:65]
  reg [63:0] counterValue; // @[BFS.scala 1120:29]
  wire  _controls_io_writeFlag_0_T = status == 3'h3; // @[BFS.scala 1123:38]
  wire  _controls_io_writeFlag_0_T_1 = status == 3'h2; // @[BFS.scala 1123:59]
  wire  _controls_io_writeFlag_0_T_3 = status == 3'h2 & io_signal_ack; // @[BFS.scala 1123:70]
  wire  _controls_io_writeFlag_0_T_5 = status == 3'h6; // @[BFS.scala 1123:108]
  wire [3:0] _controls_io_wptr_0_T_3 = _controls_io_writeFlag_0_T_1 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_0_T_4 = _controls_io_writeFlag_0_T_5 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_0_T_6 = _controls_io_wptr_0_T_3 | _controls_io_wptr_0_T_4; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_5 = _controls_io_writeFlag_0_T_1 ? new_tep[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_6 = _controls_io_writeFlag_0_T_5 ? counterValue[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [1:0] _controls_io_dataIn_0_T_7 = _controls_io_writeFlag_0_T ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_0_T_8 = _controls_io_dataIn_0_T_5 | _controls_io_dataIn_0_T_6; // @[Mux.scala 27:72]
  wire [31:0] _GEN_46 = {{30'd0}, _controls_io_dataIn_0_T_7}; // @[Mux.scala 27:72]
  wire [3:0] _controls_io_wptr_1_T_1 = _controls_io_writeFlag_0_T_1 ? 4'hd : 4'hf; // @[BFS.scala 1135:29]
  wire [31:0] _controls_io_dataIn_1_T_4 = _controls_io_writeFlag_0_T_1 ? new_tep[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _controls_io_dataIn_1_T_5 = _controls_io_writeFlag_0_T_5 ? counterValue[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1 = status == 3'h0 & start; // @[BFS.scala 1141:28]
  wire  _T_2 = status == 3'h4; // @[BFS.scala 1143:21]
  wire [2:0] _GEN_0 = io_unvisited_size == 32'h0 ? 3'h6 : 3'h1; // @[BFS.scala 1148:36 BFS.scala 1149:14 BFS.scala 1151:14]
  wire [2:0] _GEN_1 = _controls_io_writeFlag_0_T_5 ? 3'h5 : status; // @[BFS.scala 1155:40 BFS.scala 1156:12 BFS.scala 1116:23]
  wire [2:0] _GEN_2 = status == 3'h5 & io_flush_cache_end ? 3'h3 : _GEN_1; // @[BFS.scala 1153:62 BFS.scala 1154:12]
  wire [2:0] _GEN_3 = _controls_io_writeFlag_0_T_3 ? _GEN_0 : _GEN_2; // @[BFS.scala 1147:60]
  wire  _GEN_7 = io_fin_0 | FIN_0; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_9 = io_fin_1 | FIN_1; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_11 = io_fin_2 | FIN_2; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_13 = io_fin_3 | FIN_3; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_15 = io_fin_4 | FIN_4; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_17 = io_fin_5 | FIN_5; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_19 = io_fin_6 | FIN_6; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_21 = io_fin_7 | FIN_7; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_23 = io_fin_8 | FIN_8; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_25 = io_fin_9 | FIN_9; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_27 = io_fin_10 | FIN_10; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_29 = io_fin_11 | FIN_11; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_31 = io_fin_12 | FIN_12; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_33 = io_fin_13 | FIN_13; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_35 = io_fin_14 | FIN_14; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_37 = io_fin_15 | FIN_15; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire  _GEN_39 = io_fin_16 | FIN_16; // @[BFS.scala 1165:28 BFS.scala 1166:11 BFS.scala 1118:20]
  wire [31:0] _level_T_1 = level + 32'h1; // @[BFS.scala 1172:20]
  wire  global_start = _controls_io_writeFlag_0_T_3 & level == 32'hffffffff; // @[BFS.scala 1177:68]
  wire [63:0] _counterValue_T_1 = counterValue + 64'h1; // @[BFS.scala 1181:34]
  reg [63:0] performanceValue_0; // @[BFS.scala 1184:33]
  wire [63:0] _performanceValue_0_T_1 = performanceValue_0 + 64'h1; // @[BFS.scala 1191:52]
  LookupTable controls ( // @[BFS.scala 1105:24]
    .clock(controls_clock),
    .reset(controls_reset),
    .io_data_0(controls_io_data_0),
    .io_data_1(controls_io_data_1),
    .io_data_2(controls_io_data_2),
    .io_data_3(controls_io_data_3),
    .io_data_4(controls_io_data_4),
    .io_data_5(controls_io_data_5),
    .io_data_6(controls_io_data_6),
    .io_data_7(controls_io_data_7),
    .io_data_8(controls_io_data_8),
    .io_data_9(controls_io_data_9),
    .io_data_10(controls_io_data_10),
    .io_data_11(controls_io_data_11),
    .io_data_12(controls_io_data_12),
    .io_data_13(controls_io_data_13),
    .io_data_16(controls_io_data_16),
    .io_data_17(controls_io_data_17),
    .io_data_18(controls_io_data_18),
    .io_dataIn_0(controls_io_dataIn_0),
    .io_dataIn_1(controls_io_dataIn_1),
    .io_writeFlag_0(controls_io_writeFlag_0),
    .io_writeFlag_1(controls_io_writeFlag_1),
    .io_wptr_0(controls_io_wptr_0),
    .io_wptr_1(controls_io_wptr_1),
    .config_awaddr(controls_config_awaddr),
    .config_awvalid(controls_config_awvalid),
    .config_awready(controls_config_awready),
    .config_araddr(controls_config_araddr),
    .config_arvalid(controls_config_arvalid),
    .config_arready(controls_config_arready),
    .config_wdata(controls_config_wdata),
    .config_wvalid(controls_config_wvalid),
    .config_wready(controls_config_wready),
    .config_rdata(controls_config_rdata),
    .config_rvalid(controls_config_rvalid),
    .config_rready(controls_config_rready),
    .config_bvalid(controls_config_bvalid),
    .config_bready(controls_config_bready)
  );
  assign io_data_0 = controls_io_data_0; // @[BFS.scala 1197:11]
  assign io_data_1 = controls_io_data_1; // @[BFS.scala 1197:11]
  assign io_data_2 = controls_io_data_2; // @[BFS.scala 1197:11]
  assign io_data_3 = controls_io_data_3; // @[BFS.scala 1197:11]
  assign io_data_4 = controls_io_data_4; // @[BFS.scala 1197:11]
  assign io_data_5 = controls_io_data_5; // @[BFS.scala 1197:11]
  assign io_data_6 = controls_io_data_6; // @[BFS.scala 1197:11]
  assign io_data_7 = controls_io_data_7; // @[BFS.scala 1197:11]
  assign io_data_8 = controls_io_data_8; // @[BFS.scala 1197:11]
  assign io_data_9 = controls_io_data_9; // @[BFS.scala 1197:11]
  assign io_data_10 = controls_io_data_10; // @[BFS.scala 1197:11]
  assign io_data_11 = controls_io_data_11; // @[BFS.scala 1197:11]
  assign io_data_16 = controls_io_data_16; // @[BFS.scala 1197:11]
  assign io_data_17 = controls_io_data_17; // @[BFS.scala 1197:11]
  assign io_data_18 = controls_io_data_18; // @[BFS.scala 1197:11]
  assign io_signal = _T_2 | _controls_io_writeFlag_0_T_1 & io_unvisited_size != 32'h0; // @[BFS.scala 1196:36]
  assign io_start = status == 3'h4; // @[BFS.scala 1199:22]
  assign io_level = level; // @[BFS.scala 1198:12]
  assign io_config_awready = controls_config_awready; // @[BFS.scala 1122:19]
  assign io_config_arready = controls_config_arready; // @[BFS.scala 1122:19]
  assign io_config_wready = controls_config_wready; // @[BFS.scala 1122:19]
  assign io_config_rdata = controls_config_rdata; // @[BFS.scala 1122:19]
  assign io_config_rvalid = controls_config_rvalid; // @[BFS.scala 1122:19]
  assign io_config_bvalid = controls_config_bvalid; // @[BFS.scala 1122:19]
  assign io_flush_cache = status == 3'h5; // @[BFS.scala 1200:28]
  assign controls_clock = clock;
  assign controls_reset = reset;
  assign controls_io_dataIn_0 = _controls_io_dataIn_0_T_8 | _GEN_46; // @[Mux.scala 27:72]
  assign controls_io_dataIn_1 = _controls_io_dataIn_1_T_4 | _controls_io_dataIn_1_T_5; // @[Mux.scala 27:72]
  assign controls_io_writeFlag_0 = status == 3'h3 | status == 3'h2 & io_signal_ack | status == 3'h6; // @[BFS.scala 1123:99]
  assign controls_io_writeFlag_1 = _controls_io_writeFlag_0_T_3 | _controls_io_writeFlag_0_T_5; // @[BFS.scala 1134:79]
  assign controls_io_wptr_0 = {{1'd0}, _controls_io_wptr_0_T_6}; // @[Mux.scala 27:72]
  assign controls_io_wptr_1 = {{1'd0}, _controls_io_wptr_1_T_1}; // @[BFS.scala 1135:29]
  assign controls_config_awaddr = io_config_awaddr; // @[BFS.scala 1122:19]
  assign controls_config_awvalid = io_config_awvalid; // @[BFS.scala 1122:19]
  assign controls_config_araddr = io_config_araddr; // @[BFS.scala 1122:19]
  assign controls_config_arvalid = io_config_arvalid; // @[BFS.scala 1122:19]
  assign controls_config_wdata = io_config_wdata; // @[BFS.scala 1122:19]
  assign controls_config_wvalid = io_config_wvalid; // @[BFS.scala 1122:19]
  assign controls_config_rready = io_config_rready; // @[BFS.scala 1122:19]
  assign controls_config_bready = io_config_bready; // @[BFS.scala 1122:19]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 1106:22]
      level <= 32'h0; // @[BFS.scala 1106:22]
    end else if (_controls_io_writeFlag_0_T_3) begin // @[BFS.scala 1171:54]
      level <= _level_T_1; // @[BFS.scala 1172:11]
    end else if (_T_1) begin // @[BFS.scala 1173:43]
      level <= 32'hffffffff; // @[BFS.scala 1174:11]
    end
    if (reset) begin // @[BFS.scala 1116:23]
      status <= 3'h0; // @[BFS.scala 1116:23]
    end else if (status == 3'h0 & start) begin // @[BFS.scala 1141:37]
      status <= 3'h4; // @[BFS.scala 1142:12]
    end else if (status == 3'h4) begin // @[BFS.scala 1143:34]
      status <= 3'h1; // @[BFS.scala 1144:12]
    end else if (status == 3'h1 & (FIN_0 & FIN_1 & FIN_2 & FIN_3 & FIN_4 & FIN_5 & FIN_6 & FIN_7 & FIN_8 & FIN_9 &
      FIN_10 & FIN_11 & FIN_12 & FIN_13 & FIN_14 & FIN_15 & FIN_16)) begin // @[BFS.scala 1145:51]
      status <= 3'h2; // @[BFS.scala 1146:12]
    end else begin
      status <= _GEN_3;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_0 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_0 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_0 <= _GEN_7;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_1 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_1 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_1 <= _GEN_9;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_2 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_2 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_2 <= _GEN_11;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_3 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_3 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_3 <= _GEN_13;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_4 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_4 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_4 <= _GEN_15;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_5 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_5 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_5 <= _GEN_17;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_6 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_6 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_6 <= _GEN_19;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_7 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_7 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_7 <= _GEN_21;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_8 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_8 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_8 <= _GEN_23;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_9 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_9 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_9 <= _GEN_25;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_10 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_10 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_10 <= _GEN_27;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_11 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_11 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_11 <= _GEN_29;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_12 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_12 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_12 <= _GEN_31;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_13 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_13 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_13 <= _GEN_33;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_14 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_14 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_14 <= _GEN_35;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_15 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_15 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_15 <= _GEN_37;
    end
    if (reset) begin // @[BFS.scala 1118:20]
      FIN_16 <= 1'h0; // @[BFS.scala 1118:20]
    end else if (io_signal) begin // @[BFS.scala 1163:22]
      FIN_16 <= 1'h0; // @[BFS.scala 1164:11]
    end else begin
      FIN_16 <= _GEN_39;
    end
    if (reset) begin // @[BFS.scala 1120:29]
      counterValue <= 64'h0; // @[BFS.scala 1120:29]
    end else if (global_start) begin // @[BFS.scala 1178:22]
      counterValue <= 64'h0; // @[BFS.scala 1179:18]
    end else begin
      counterValue <= _counterValue_T_1; // @[BFS.scala 1181:18]
    end
    if (reset) begin // @[BFS.scala 1184:33]
      performanceValue_0 <= 64'h0; // @[BFS.scala 1184:33]
    end else if (global_start) begin // @[BFS.scala 1188:26]
      performanceValue_0 <= 64'h0; // @[BFS.scala 1189:29]
    end else if (io_performance_0) begin // @[BFS.scala 1190:20]
      performanceValue_0 <= _performanceValue_0_T_1; // @[BFS.scala 1191:29]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  level = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  status = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  FIN_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  FIN_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  FIN_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  FIN_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  FIN_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  FIN_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  FIN_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  FIN_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  FIN_8 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  FIN_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  FIN_10 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  FIN_11 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  FIN_12 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  FIN_13 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  FIN_14 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  FIN_15 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  FIN_16 = _RAND_18[0:0];
  _RAND_19 = {2{`RANDOM}};
  counterValue = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  performanceValue_0 = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pipeline(
  input         clock,
  input         reset,
  input         io_dout_ready,
  output        io_dout_valid,
  output [31:0] io_dout_bits_tdata,
  output        io_din_ready,
  input         io_din_valid,
  input  [31:0] io_din_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] data_tdata; // @[util.scala 238:21]
  reg  valid; // @[util.scala 239:22]
  reg  ready; // @[util.scala 240:22]
  reg [31:0] data2_tdata; // @[util.scala 241:22]
  reg  valid2; // @[util.scala 242:23]
  wire  _GEN_3 = ready & io_din_valid; // @[util.scala 247:22 util.scala 249:13 util.scala 252:13]
  assign io_dout_valid = valid; // @[util.scala 268:17]
  assign io_dout_bits_tdata = data_tdata; // @[util.scala 269:16]
  assign io_din_ready = ready; // @[util.scala 267:16]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 238:21]
      data_tdata <= 32'h0; // @[util.scala 238:21]
    end else if (io_dout_ready) begin // @[util.scala 243:22]
      if (valid2) begin // @[util.scala 244:17]
        data_tdata <= data2_tdata; // @[util.scala 245:12]
      end else if (ready) begin // @[util.scala 247:22]
        data_tdata <= io_din_bits_tdata; // @[util.scala 248:12]
      end else begin
        data_tdata <= 32'h0; // @[util.scala 251:12]
      end
    end
    if (reset) begin // @[util.scala 239:22]
      valid <= 1'h0; // @[util.scala 239:22]
    end else if (io_dout_ready) begin // @[util.scala 243:22]
      if (valid2) begin // @[util.scala 244:17]
        valid <= valid2; // @[util.scala 246:13]
      end else begin
        valid <= _GEN_3;
      end
    end
    if (reset) begin // @[util.scala 240:22]
      ready <= 1'h0; // @[util.scala 240:22]
    end else begin
      ready <= io_dout_ready; // @[util.scala 255:9]
    end
    if (reset) begin // @[util.scala 241:22]
      data2_tdata <= 32'h0; // @[util.scala 241:22]
    end else if (~io_dout_ready & ready) begin // @[util.scala 258:33]
      data2_tdata <= io_din_bits_tdata; // @[util.scala 259:11]
    end else if (io_dout_ready) begin // @[util.scala 261:28]
      data2_tdata <= 32'h0; // @[util.scala 263:11]
    end
    if (reset) begin // @[util.scala 242:23]
      valid2 <= 1'h0; // @[util.scala 242:23]
    end else if (~io_dout_ready & ready) begin // @[util.scala 258:33]
      valid2 <= io_din_valid; // @[util.scala 260:12]
    end else if (io_dout_ready) begin // @[util.scala 261:28]
      valid2 <= 1'h0; // @[util.scala 264:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_tdata = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ready = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  data2_tdata = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  valid2 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multi_channel_fifo(
  input          clock,
  input          reset,
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [31:0]  io_in_0_bits_tdata,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [31:0]  io_in_1_bits_tdata,
  output         io_in_2_ready,
  input          io_in_2_valid,
  input  [31:0]  io_in_2_bits_tdata,
  output         io_in_3_ready,
  input          io_in_3_valid,
  input  [31:0]  io_in_3_bits_tdata,
  output         io_in_4_ready,
  input          io_in_4_valid,
  input  [31:0]  io_in_4_bits_tdata,
  output         io_in_5_ready,
  input          io_in_5_valid,
  input  [31:0]  io_in_5_bits_tdata,
  output         io_in_6_ready,
  input          io_in_6_valid,
  input  [31:0]  io_in_6_bits_tdata,
  output         io_in_7_ready,
  input          io_in_7_valid,
  input  [31:0]  io_in_7_bits_tdata,
  output         io_in_8_ready,
  input          io_in_8_valid,
  input  [31:0]  io_in_8_bits_tdata,
  output         io_in_9_ready,
  input          io_in_9_valid,
  input  [31:0]  io_in_9_bits_tdata,
  output         io_in_10_ready,
  input          io_in_10_valid,
  input  [31:0]  io_in_10_bits_tdata,
  output         io_in_11_ready,
  input          io_in_11_valid,
  input  [31:0]  io_in_11_bits_tdata,
  output         io_in_12_ready,
  input          io_in_12_valid,
  input  [31:0]  io_in_12_bits_tdata,
  output         io_in_13_ready,
  input          io_in_13_valid,
  input  [31:0]  io_in_13_bits_tdata,
  output         io_in_14_ready,
  input          io_in_14_valid,
  input  [31:0]  io_in_14_bits_tdata,
  output         io_in_15_ready,
  input          io_in_15_valid,
  input  [31:0]  io_in_15_bits_tdata,
  output         io_out_full,
  input  [511:0] io_out_din,
  input          io_out_wr_en,
  output [511:0] io_out_dout,
  input          io_out_rd_en,
  output [8:0]   io_out_data_count,
  output         io_out_valid,
  input          io_flush,
  input          io_is_current_tier
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  collector_fifos_0_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_0_din; // @[BFS.scala 826:16]
  wire  collector_fifos_0_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_0_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_0_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_0_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_0_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_0_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_0_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_0_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_1_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_1_din; // @[BFS.scala 826:16]
  wire  collector_fifos_1_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_1_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_1_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_1_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_1_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_1_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_1_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_1_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_2_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_2_din; // @[BFS.scala 826:16]
  wire  collector_fifos_2_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_2_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_2_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_2_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_2_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_2_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_2_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_2_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_3_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_3_din; // @[BFS.scala 826:16]
  wire  collector_fifos_3_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_3_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_3_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_3_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_3_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_3_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_3_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_3_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_4_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_4_din; // @[BFS.scala 826:16]
  wire  collector_fifos_4_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_4_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_4_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_4_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_4_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_4_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_4_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_4_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_5_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_5_din; // @[BFS.scala 826:16]
  wire  collector_fifos_5_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_5_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_5_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_5_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_5_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_5_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_5_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_5_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_6_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_6_din; // @[BFS.scala 826:16]
  wire  collector_fifos_6_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_6_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_6_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_6_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_6_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_6_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_6_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_6_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_7_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_7_din; // @[BFS.scala 826:16]
  wire  collector_fifos_7_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_7_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_7_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_7_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_7_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_7_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_7_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_7_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_8_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_8_din; // @[BFS.scala 826:16]
  wire  collector_fifos_8_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_8_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_8_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_8_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_8_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_8_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_8_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_8_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_9_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_9_din; // @[BFS.scala 826:16]
  wire  collector_fifos_9_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_9_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_9_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_9_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_9_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_9_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_9_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_9_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_10_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_10_din; // @[BFS.scala 826:16]
  wire  collector_fifos_10_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_10_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_10_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_10_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_10_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_10_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_10_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_10_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_11_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_11_din; // @[BFS.scala 826:16]
  wire  collector_fifos_11_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_11_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_11_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_11_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_11_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_11_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_11_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_11_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_12_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_12_din; // @[BFS.scala 826:16]
  wire  collector_fifos_12_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_12_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_12_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_12_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_12_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_12_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_12_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_12_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_13_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_13_din; // @[BFS.scala 826:16]
  wire  collector_fifos_13_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_13_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_13_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_13_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_13_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_13_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_13_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_13_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_14_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_14_din; // @[BFS.scala 826:16]
  wire  collector_fifos_14_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_14_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_14_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_14_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_14_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_14_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_14_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_14_valid; // @[BFS.scala 826:16]
  wire  collector_fifos_15_full; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_15_din; // @[BFS.scala 826:16]
  wire  collector_fifos_15_wr_en; // @[BFS.scala 826:16]
  wire  collector_fifos_15_empty; // @[BFS.scala 826:16]
  wire [31:0] collector_fifos_15_dout; // @[BFS.scala 826:16]
  wire  collector_fifos_15_rd_en; // @[BFS.scala 826:16]
  wire [4:0] collector_fifos_15_data_count; // @[BFS.scala 826:16]
  wire  collector_fifos_15_clk; // @[BFS.scala 826:16]
  wire  collector_fifos_15_srst; // @[BFS.scala 826:16]
  wire  collector_fifos_15_valid; // @[BFS.scala 826:16]
  wire  in_pipeline_0_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_0_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_0_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_0_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_0_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_0_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_0_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_0_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_1_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_1_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_1_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_1_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_1_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_1_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_1_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_1_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_2_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_2_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_2_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_2_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_2_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_2_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_2_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_2_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_3_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_3_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_3_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_3_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_3_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_3_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_3_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_3_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_4_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_4_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_4_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_4_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_4_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_4_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_4_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_4_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_5_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_5_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_5_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_5_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_5_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_5_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_5_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_5_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_6_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_6_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_6_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_6_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_6_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_6_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_6_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_6_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_7_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_7_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_7_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_7_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_7_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_7_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_7_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_7_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_8_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_8_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_8_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_8_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_8_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_8_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_8_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_8_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_9_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_9_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_9_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_9_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_9_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_9_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_9_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_9_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_10_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_10_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_10_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_10_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_10_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_10_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_10_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_10_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_11_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_11_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_11_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_11_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_11_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_11_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_11_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_11_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_12_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_12_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_12_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_12_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_12_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_12_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_12_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_12_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_13_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_13_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_13_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_13_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_13_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_13_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_13_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_13_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_14_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_14_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_14_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_14_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_14_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_14_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_14_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_14_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_15_clock; // @[BFS.scala 832:11]
  wire  in_pipeline_15_reset; // @[BFS.scala 832:11]
  wire  in_pipeline_15_io_dout_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_15_io_dout_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_15_io_dout_bits_tdata; // @[BFS.scala 832:11]
  wire  in_pipeline_15_io_din_ready; // @[BFS.scala 832:11]
  wire  in_pipeline_15_io_din_valid; // @[BFS.scala 832:11]
  wire [31:0] in_pipeline_15_io_din_bits_tdata; // @[BFS.scala 832:11]
  wire  _fifos_ready_T_15 = ~collector_fifos_15_full; // @[BFS.scala 828:70]
  wire  fifos_ready = ~collector_fifos_0_full & ~collector_fifos_1_full & ~collector_fifos_2_full & ~
    collector_fifos_3_full & ~collector_fifos_4_full & ~collector_fifos_5_full & ~collector_fifos_6_full & ~
    collector_fifos_7_full & ~collector_fifos_8_full & ~collector_fifos_9_full & ~collector_fifos_10_full & ~
    collector_fifos_11_full & ~collector_fifos_12_full & ~collector_fifos_13_full & ~collector_fifos_14_full &
    _fifos_ready_T_15; // @[BFS.scala 828:91]
  reg [3:0] counter; // @[BFS.scala 829:24]
  wire  _steps_T = in_pipeline_0_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire  _steps_T_2 = in_pipeline_1_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE = {{4'd0}, _steps_T}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] _steps_WIRE_1 = {{4'd0}, _steps_T_2}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_1 = _steps_WIRE + _steps_WIRE_1; // @[BFS.scala 842:107]
  wire  _steps_T_6 = in_pipeline_2_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_4 = {{4'd0}, _steps_T_6}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_2 = steps_1 + _steps_WIRE_4; // @[BFS.scala 842:107]
  wire  _steps_T_13 = in_pipeline_3_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_8 = {{4'd0}, _steps_T_13}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_3 = steps_2 + _steps_WIRE_8; // @[BFS.scala 842:107]
  wire  _steps_T_23 = in_pipeline_4_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_13 = {{4'd0}, _steps_T_23}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_4 = steps_3 + _steps_WIRE_13; // @[BFS.scala 842:107]
  wire  _steps_T_36 = in_pipeline_5_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_19 = {{4'd0}, _steps_T_36}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_5 = steps_4 + _steps_WIRE_19; // @[BFS.scala 842:107]
  wire  _steps_T_52 = in_pipeline_6_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_26 = {{4'd0}, _steps_T_52}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_6 = steps_5 + _steps_WIRE_26; // @[BFS.scala 842:107]
  wire  _steps_T_71 = in_pipeline_7_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_34 = {{4'd0}, _steps_T_71}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_7 = steps_6 + _steps_WIRE_34; // @[BFS.scala 842:107]
  wire  _steps_T_93 = in_pipeline_8_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_43 = {{4'd0}, _steps_T_93}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_8 = steps_7 + _steps_WIRE_43; // @[BFS.scala 842:107]
  wire  _steps_T_118 = in_pipeline_9_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_53 = {{4'd0}, _steps_T_118}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_9 = steps_8 + _steps_WIRE_53; // @[BFS.scala 842:107]
  wire  _steps_T_146 = in_pipeline_10_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_64 = {{4'd0}, _steps_T_146}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_10 = steps_9 + _steps_WIRE_64; // @[BFS.scala 842:107]
  wire  _steps_T_177 = in_pipeline_11_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_76 = {{4'd0}, _steps_T_177}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_11 = steps_10 + _steps_WIRE_76; // @[BFS.scala 842:107]
  wire  _steps_T_211 = in_pipeline_12_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_89 = {{4'd0}, _steps_T_211}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_12 = steps_11 + _steps_WIRE_89; // @[BFS.scala 842:107]
  wire  _steps_T_248 = in_pipeline_13_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_103 = {{4'd0}, _steps_T_248}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_13 = steps_12 + _steps_WIRE_103; // @[BFS.scala 842:107]
  wire  _steps_T_288 = in_pipeline_14_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_118 = {{4'd0}, _steps_T_288}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_14 = steps_13 + _steps_WIRE_118; // @[BFS.scala 842:107]
  wire  _steps_T_331 = in_pipeline_15_io_dout_valid & fifos_ready; // @[BFS.scala 842:62]
  wire [4:0] _steps_WIRE_134 = {{4'd0}, _steps_T_331}; // @[BFS.scala 842:86 BFS.scala 842:86]
  wire [4:0] steps_15 = steps_14 + _steps_WIRE_134; // @[BFS.scala 842:107]
  wire [4:0] _GEN_2 = {{1'd0}, counter}; // @[BFS.scala 847:15]
  wire [4:0] _counter_T_1 = _GEN_2 + steps_15; // @[BFS.scala 847:15]
  wire [4:0] _counter_T_6 = _counter_T_1 - 5'h10; // @[BFS.scala 847:44]
  wire [4:0] _counter_T_9 = _counter_T_1 >= 5'h10 ? _counter_T_6 : _counter_T_1; // @[BFS.scala 847:8]
  wire [3:0] _GEN_0 = io_flush ? 4'h0 : counter; // @[BFS.scala 855:23 BFS.scala 856:13 BFS.scala 829:24]
  wire [4:0] _GEN_1 = steps_15 != 5'h0 ? _counter_T_9 : {{1'd0}, _GEN_0}; // @[BFS.scala 853:39 BFS.scala 854:13]
  wire [3:0] _fifo_in_data_T_2 = 4'h0 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_4 = 5'h10 - _GEN_2; // @[BFS.scala 850:49]
  wire [5:0] _fifo_in_data_T_5 = {{1'd0}, _fifo_in_data_T_4}; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_7 = counter <= 4'h0 ? {{1'd0}, _fifo_in_data_T_2} : _fifo_in_data_T_5[4:0]; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_9 = _fifo_in_data_T_7 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_10 = _fifo_in_data_T_9 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_21 = _fifo_in_data_T_9 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_32 = _fifo_in_data_T_9 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_43 = _fifo_in_data_T_9 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_54 = _fifo_in_data_T_9 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_65 = _fifo_in_data_T_9 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_76 = _fifo_in_data_T_9 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_87 = _fifo_in_data_T_9 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_98 = _fifo_in_data_T_9 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_109 = _fifo_in_data_T_9 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_120 = _fifo_in_data_T_9 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_131 = _fifo_in_data_T_9 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_142 = _fifo_in_data_T_9 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_153 = _fifo_in_data_T_9 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_164 = _fifo_in_data_T_9 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_175 = _fifo_in_data_T_9 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_176 = _fifo_in_data_T_175 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_177 = _fifo_in_data_T_164 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_176; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_178 = _fifo_in_data_T_153 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_177; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_179 = _fifo_in_data_T_142 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_178; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_180 = _fifo_in_data_T_131 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_179; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_181 = _fifo_in_data_T_120 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_180; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_182 = _fifo_in_data_T_109 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_181; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_183 = _fifo_in_data_T_98 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_182; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_184 = _fifo_in_data_T_87 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_183; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_185 = _fifo_in_data_T_76 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_184; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_186 = _fifo_in_data_T_65 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_185; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_187 = _fifo_in_data_T_54 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_186; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_188 = _fifo_in_data_T_43 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_187; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_189 = _fifo_in_data_T_32 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_188; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_190 = _fifo_in_data_T_21 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_189; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data = _fifo_in_data_T_10 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_190; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_177 = _fifo_in_data_T_164 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_175 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_178 = _fifo_in_data_T_153 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_177; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_179 = _fifo_in_data_T_142 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_178; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_180 = _fifo_in_data_T_131 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_179; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_181 = _fifo_in_data_T_120 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_180; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_182 = _fifo_in_data_T_109 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_181; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_183 = _fifo_in_data_T_98 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_182; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_184 = _fifo_in_data_T_87 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_183; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_185 = _fifo_in_data_T_76 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_184; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_186 = _fifo_in_data_T_65 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_185; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_187 = _fifo_in_data_T_54 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_186; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_188 = _fifo_in_data_T_43 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_187; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_189 = _fifo_in_data_T_32 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_188; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_190 = _fifo_in_data_T_21 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_189; // @[Mux.scala 98:16]
  wire  fifo_in_valid = _fifo_in_data_T_10 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_190; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_193 = 4'h1 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_197 = _fifo_in_data_T_4 + 5'h1; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_198 = counter <= 4'h1 ? {{1'd0}, _fifo_in_data_T_193} : _fifo_in_data_T_197; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_200 = _fifo_in_data_T_198 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_201 = _fifo_in_data_T_200 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_212 = _fifo_in_data_T_200 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_223 = _fifo_in_data_T_200 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_234 = _fifo_in_data_T_200 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_245 = _fifo_in_data_T_200 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_256 = _fifo_in_data_T_200 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_267 = _fifo_in_data_T_200 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_278 = _fifo_in_data_T_200 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_289 = _fifo_in_data_T_200 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_300 = _fifo_in_data_T_200 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_311 = _fifo_in_data_T_200 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_322 = _fifo_in_data_T_200 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_333 = _fifo_in_data_T_200 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_344 = _fifo_in_data_T_200 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_355 = _fifo_in_data_T_200 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_366 = _fifo_in_data_T_200 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_367 = _fifo_in_data_T_366 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_368 = _fifo_in_data_T_355 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_367; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_369 = _fifo_in_data_T_344 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_368; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_370 = _fifo_in_data_T_333 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_369; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_371 = _fifo_in_data_T_322 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_370; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_372 = _fifo_in_data_T_311 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_371; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_373 = _fifo_in_data_T_300 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_372; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_374 = _fifo_in_data_T_289 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_373; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_375 = _fifo_in_data_T_278 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_374; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_376 = _fifo_in_data_T_267 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_375; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_377 = _fifo_in_data_T_256 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_376; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_378 = _fifo_in_data_T_245 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_377; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_379 = _fifo_in_data_T_234 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_378; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_380 = _fifo_in_data_T_223 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_379; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_381 = _fifo_in_data_T_212 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_380; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_1 = _fifo_in_data_T_201 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_381; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_368 = _fifo_in_data_T_355 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_366 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_369 = _fifo_in_data_T_344 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_368; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_370 = _fifo_in_data_T_333 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_369; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_371 = _fifo_in_data_T_322 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_370; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_372 = _fifo_in_data_T_311 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_371; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_373 = _fifo_in_data_T_300 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_372; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_374 = _fifo_in_data_T_289 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_373; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_375 = _fifo_in_data_T_278 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_374; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_376 = _fifo_in_data_T_267 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_375; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_377 = _fifo_in_data_T_256 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_376; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_378 = _fifo_in_data_T_245 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_377; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_379 = _fifo_in_data_T_234 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_378; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_380 = _fifo_in_data_T_223 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_379; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_381 = _fifo_in_data_T_212 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_380; // @[Mux.scala 98:16]
  wire  fifo_in_valid_1 = _fifo_in_data_T_201 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_381; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_384 = 4'h2 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_388 = _fifo_in_data_T_4 + 5'h2; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_389 = counter <= 4'h2 ? {{1'd0}, _fifo_in_data_T_384} : _fifo_in_data_T_388; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_391 = _fifo_in_data_T_389 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_392 = _fifo_in_data_T_391 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_403 = _fifo_in_data_T_391 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_414 = _fifo_in_data_T_391 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_425 = _fifo_in_data_T_391 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_436 = _fifo_in_data_T_391 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_447 = _fifo_in_data_T_391 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_458 = _fifo_in_data_T_391 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_469 = _fifo_in_data_T_391 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_480 = _fifo_in_data_T_391 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_491 = _fifo_in_data_T_391 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_502 = _fifo_in_data_T_391 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_513 = _fifo_in_data_T_391 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_524 = _fifo_in_data_T_391 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_535 = _fifo_in_data_T_391 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_546 = _fifo_in_data_T_391 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_557 = _fifo_in_data_T_391 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_558 = _fifo_in_data_T_557 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_559 = _fifo_in_data_T_546 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_558; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_560 = _fifo_in_data_T_535 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_559; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_561 = _fifo_in_data_T_524 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_560; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_562 = _fifo_in_data_T_513 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_561; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_563 = _fifo_in_data_T_502 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_562; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_564 = _fifo_in_data_T_491 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_563; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_565 = _fifo_in_data_T_480 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_564; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_566 = _fifo_in_data_T_469 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_565; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_567 = _fifo_in_data_T_458 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_566; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_568 = _fifo_in_data_T_447 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_567; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_569 = _fifo_in_data_T_436 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_568; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_570 = _fifo_in_data_T_425 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_569; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_571 = _fifo_in_data_T_414 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_570; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_572 = _fifo_in_data_T_403 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_571; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_2 = _fifo_in_data_T_392 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_572; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_559 = _fifo_in_data_T_546 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_557 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_560 = _fifo_in_data_T_535 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_559; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_561 = _fifo_in_data_T_524 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_560; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_562 = _fifo_in_data_T_513 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_561; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_563 = _fifo_in_data_T_502 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_562; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_564 = _fifo_in_data_T_491 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_563; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_565 = _fifo_in_data_T_480 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_564; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_566 = _fifo_in_data_T_469 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_565; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_567 = _fifo_in_data_T_458 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_566; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_568 = _fifo_in_data_T_447 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_567; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_569 = _fifo_in_data_T_436 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_568; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_570 = _fifo_in_data_T_425 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_569; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_571 = _fifo_in_data_T_414 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_570; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_572 = _fifo_in_data_T_403 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_571; // @[Mux.scala 98:16]
  wire  fifo_in_valid_2 = _fifo_in_data_T_392 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_572; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_575 = 4'h3 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_579 = _fifo_in_data_T_4 + 5'h3; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_580 = counter <= 4'h3 ? {{1'd0}, _fifo_in_data_T_575} : _fifo_in_data_T_579; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_582 = _fifo_in_data_T_580 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_583 = _fifo_in_data_T_582 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_594 = _fifo_in_data_T_582 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_605 = _fifo_in_data_T_582 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_616 = _fifo_in_data_T_582 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_627 = _fifo_in_data_T_582 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_638 = _fifo_in_data_T_582 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_649 = _fifo_in_data_T_582 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_660 = _fifo_in_data_T_582 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_671 = _fifo_in_data_T_582 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_682 = _fifo_in_data_T_582 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_693 = _fifo_in_data_T_582 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_704 = _fifo_in_data_T_582 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_715 = _fifo_in_data_T_582 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_726 = _fifo_in_data_T_582 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_737 = _fifo_in_data_T_582 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_748 = _fifo_in_data_T_582 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_749 = _fifo_in_data_T_748 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_750 = _fifo_in_data_T_737 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_749; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_751 = _fifo_in_data_T_726 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_750; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_752 = _fifo_in_data_T_715 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_751; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_753 = _fifo_in_data_T_704 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_752; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_754 = _fifo_in_data_T_693 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_753; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_755 = _fifo_in_data_T_682 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_754; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_756 = _fifo_in_data_T_671 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_755; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_757 = _fifo_in_data_T_660 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_756; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_758 = _fifo_in_data_T_649 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_757; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_759 = _fifo_in_data_T_638 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_758; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_760 = _fifo_in_data_T_627 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_759; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_761 = _fifo_in_data_T_616 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_760; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_762 = _fifo_in_data_T_605 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_761; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_763 = _fifo_in_data_T_594 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_762; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_3 = _fifo_in_data_T_583 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_763; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_750 = _fifo_in_data_T_737 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_748 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_751 = _fifo_in_data_T_726 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_750; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_752 = _fifo_in_data_T_715 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_751; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_753 = _fifo_in_data_T_704 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_752; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_754 = _fifo_in_data_T_693 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_753; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_755 = _fifo_in_data_T_682 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_754; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_756 = _fifo_in_data_T_671 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_755; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_757 = _fifo_in_data_T_660 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_756; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_758 = _fifo_in_data_T_649 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_757; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_759 = _fifo_in_data_T_638 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_758; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_760 = _fifo_in_data_T_627 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_759; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_761 = _fifo_in_data_T_616 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_760; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_762 = _fifo_in_data_T_605 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_761; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_763 = _fifo_in_data_T_594 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_762; // @[Mux.scala 98:16]
  wire  fifo_in_valid_3 = _fifo_in_data_T_583 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_763; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_766 = 4'h4 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_770 = _fifo_in_data_T_4 + 5'h4; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_771 = counter <= 4'h4 ? {{1'd0}, _fifo_in_data_T_766} : _fifo_in_data_T_770; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_773 = _fifo_in_data_T_771 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_774 = _fifo_in_data_T_773 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_785 = _fifo_in_data_T_773 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_796 = _fifo_in_data_T_773 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_807 = _fifo_in_data_T_773 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_818 = _fifo_in_data_T_773 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_829 = _fifo_in_data_T_773 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_840 = _fifo_in_data_T_773 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_851 = _fifo_in_data_T_773 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_862 = _fifo_in_data_T_773 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_873 = _fifo_in_data_T_773 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_884 = _fifo_in_data_T_773 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_895 = _fifo_in_data_T_773 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_906 = _fifo_in_data_T_773 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_917 = _fifo_in_data_T_773 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_928 = _fifo_in_data_T_773 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_939 = _fifo_in_data_T_773 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_940 = _fifo_in_data_T_939 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_941 = _fifo_in_data_T_928 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_940; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_942 = _fifo_in_data_T_917 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_941; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_943 = _fifo_in_data_T_906 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_942; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_944 = _fifo_in_data_T_895 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_943; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_945 = _fifo_in_data_T_884 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_944; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_946 = _fifo_in_data_T_873 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_945; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_947 = _fifo_in_data_T_862 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_946; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_948 = _fifo_in_data_T_851 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_947; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_949 = _fifo_in_data_T_840 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_948; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_950 = _fifo_in_data_T_829 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_949; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_951 = _fifo_in_data_T_818 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_950; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_952 = _fifo_in_data_T_807 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_951; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_953 = _fifo_in_data_T_796 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_952; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_954 = _fifo_in_data_T_785 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_953; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_4 = _fifo_in_data_T_774 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_954; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_941 = _fifo_in_data_T_928 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_939 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_942 = _fifo_in_data_T_917 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_941; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_943 = _fifo_in_data_T_906 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_942; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_944 = _fifo_in_data_T_895 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_943; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_945 = _fifo_in_data_T_884 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_944; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_946 = _fifo_in_data_T_873 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_945; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_947 = _fifo_in_data_T_862 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_946; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_948 = _fifo_in_data_T_851 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_947; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_949 = _fifo_in_data_T_840 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_948; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_950 = _fifo_in_data_T_829 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_949; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_951 = _fifo_in_data_T_818 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_950; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_952 = _fifo_in_data_T_807 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_951; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_953 = _fifo_in_data_T_796 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_952; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_954 = _fifo_in_data_T_785 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_953; // @[Mux.scala 98:16]
  wire  fifo_in_valid_4 = _fifo_in_data_T_774 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_954; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_957 = 4'h5 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_961 = _fifo_in_data_T_4 + 5'h5; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_962 = counter <= 4'h5 ? {{1'd0}, _fifo_in_data_T_957} : _fifo_in_data_T_961; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_964 = _fifo_in_data_T_962 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_965 = _fifo_in_data_T_964 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_976 = _fifo_in_data_T_964 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_987 = _fifo_in_data_T_964 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_998 = _fifo_in_data_T_964 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1009 = _fifo_in_data_T_964 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1020 = _fifo_in_data_T_964 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1031 = _fifo_in_data_T_964 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1042 = _fifo_in_data_T_964 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1053 = _fifo_in_data_T_964 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1064 = _fifo_in_data_T_964 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1075 = _fifo_in_data_T_964 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1086 = _fifo_in_data_T_964 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1097 = _fifo_in_data_T_964 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1108 = _fifo_in_data_T_964 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1119 = _fifo_in_data_T_964 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1130 = _fifo_in_data_T_964 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1131 = _fifo_in_data_T_1130 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1132 = _fifo_in_data_T_1119 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1131; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1133 = _fifo_in_data_T_1108 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1132; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1134 = _fifo_in_data_T_1097 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1133; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1135 = _fifo_in_data_T_1086 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1134; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1136 = _fifo_in_data_T_1075 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1135; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1137 = _fifo_in_data_T_1064 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1136; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1138 = _fifo_in_data_T_1053 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1137; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1139 = _fifo_in_data_T_1042 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1138; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1140 = _fifo_in_data_T_1031 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1139; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1141 = _fifo_in_data_T_1020 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1140; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1142 = _fifo_in_data_T_1009 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1141; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1143 = _fifo_in_data_T_998 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1142; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1144 = _fifo_in_data_T_987 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1143; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1145 = _fifo_in_data_T_976 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1144; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_5 = _fifo_in_data_T_965 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1145; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1132 = _fifo_in_data_T_1119 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1130 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1133 = _fifo_in_data_T_1108 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1132; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1134 = _fifo_in_data_T_1097 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1133; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1135 = _fifo_in_data_T_1086 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1134; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1136 = _fifo_in_data_T_1075 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1135; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1137 = _fifo_in_data_T_1064 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1136; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1138 = _fifo_in_data_T_1053 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1137; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1139 = _fifo_in_data_T_1042 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1138; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1140 = _fifo_in_data_T_1031 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1139; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1141 = _fifo_in_data_T_1020 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1140; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1142 = _fifo_in_data_T_1009 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1141; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1143 = _fifo_in_data_T_998 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1142; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1144 = _fifo_in_data_T_987 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1143; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1145 = _fifo_in_data_T_976 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1144; // @[Mux.scala 98:16]
  wire  fifo_in_valid_5 = _fifo_in_data_T_965 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1145; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1148 = 4'h6 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1152 = _fifo_in_data_T_4 + 5'h6; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1153 = counter <= 4'h6 ? {{1'd0}, _fifo_in_data_T_1148} : _fifo_in_data_T_1152; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1155 = _fifo_in_data_T_1153 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1156 = _fifo_in_data_T_1155 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1167 = _fifo_in_data_T_1155 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1178 = _fifo_in_data_T_1155 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1189 = _fifo_in_data_T_1155 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1200 = _fifo_in_data_T_1155 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1211 = _fifo_in_data_T_1155 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1222 = _fifo_in_data_T_1155 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1233 = _fifo_in_data_T_1155 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1244 = _fifo_in_data_T_1155 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1255 = _fifo_in_data_T_1155 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1266 = _fifo_in_data_T_1155 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1277 = _fifo_in_data_T_1155 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1288 = _fifo_in_data_T_1155 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1299 = _fifo_in_data_T_1155 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1310 = _fifo_in_data_T_1155 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1321 = _fifo_in_data_T_1155 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1322 = _fifo_in_data_T_1321 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1323 = _fifo_in_data_T_1310 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1322; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1324 = _fifo_in_data_T_1299 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1323; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1325 = _fifo_in_data_T_1288 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1324; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1326 = _fifo_in_data_T_1277 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1325; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1327 = _fifo_in_data_T_1266 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1326; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1328 = _fifo_in_data_T_1255 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1327; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1329 = _fifo_in_data_T_1244 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1328; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1330 = _fifo_in_data_T_1233 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1329; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1331 = _fifo_in_data_T_1222 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1330; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1332 = _fifo_in_data_T_1211 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1331; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1333 = _fifo_in_data_T_1200 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1332; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1334 = _fifo_in_data_T_1189 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1333; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1335 = _fifo_in_data_T_1178 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1334; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1336 = _fifo_in_data_T_1167 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1335; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_6 = _fifo_in_data_T_1156 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1336; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1323 = _fifo_in_data_T_1310 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1321 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1324 = _fifo_in_data_T_1299 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1323; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1325 = _fifo_in_data_T_1288 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1324; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1326 = _fifo_in_data_T_1277 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1325; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1327 = _fifo_in_data_T_1266 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1326; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1328 = _fifo_in_data_T_1255 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1327; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1329 = _fifo_in_data_T_1244 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1328; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1330 = _fifo_in_data_T_1233 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1329; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1331 = _fifo_in_data_T_1222 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1330; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1332 = _fifo_in_data_T_1211 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1331; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1333 = _fifo_in_data_T_1200 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1332; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1334 = _fifo_in_data_T_1189 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1333; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1335 = _fifo_in_data_T_1178 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1334; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1336 = _fifo_in_data_T_1167 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1335; // @[Mux.scala 98:16]
  wire  fifo_in_valid_6 = _fifo_in_data_T_1156 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1336; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1339 = 4'h7 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1343 = _fifo_in_data_T_4 + 5'h7; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1344 = counter <= 4'h7 ? {{1'd0}, _fifo_in_data_T_1339} : _fifo_in_data_T_1343; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1346 = _fifo_in_data_T_1344 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1347 = _fifo_in_data_T_1346 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1358 = _fifo_in_data_T_1346 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1369 = _fifo_in_data_T_1346 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1380 = _fifo_in_data_T_1346 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1391 = _fifo_in_data_T_1346 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1402 = _fifo_in_data_T_1346 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1413 = _fifo_in_data_T_1346 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1424 = _fifo_in_data_T_1346 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1435 = _fifo_in_data_T_1346 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1446 = _fifo_in_data_T_1346 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1457 = _fifo_in_data_T_1346 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1468 = _fifo_in_data_T_1346 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1479 = _fifo_in_data_T_1346 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1490 = _fifo_in_data_T_1346 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1501 = _fifo_in_data_T_1346 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1512 = _fifo_in_data_T_1346 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1513 = _fifo_in_data_T_1512 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1514 = _fifo_in_data_T_1501 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1513; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1515 = _fifo_in_data_T_1490 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1514; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1516 = _fifo_in_data_T_1479 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1515; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1517 = _fifo_in_data_T_1468 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1516; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1518 = _fifo_in_data_T_1457 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1517; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1519 = _fifo_in_data_T_1446 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1518; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1520 = _fifo_in_data_T_1435 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1519; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1521 = _fifo_in_data_T_1424 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1520; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1522 = _fifo_in_data_T_1413 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1521; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1523 = _fifo_in_data_T_1402 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1522; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1524 = _fifo_in_data_T_1391 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1523; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1525 = _fifo_in_data_T_1380 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1524; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1526 = _fifo_in_data_T_1369 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1525; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1527 = _fifo_in_data_T_1358 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1526; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_7 = _fifo_in_data_T_1347 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1527; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1514 = _fifo_in_data_T_1501 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1512 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1515 = _fifo_in_data_T_1490 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1514; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1516 = _fifo_in_data_T_1479 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1515; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1517 = _fifo_in_data_T_1468 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1516; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1518 = _fifo_in_data_T_1457 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1517; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1519 = _fifo_in_data_T_1446 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1518; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1520 = _fifo_in_data_T_1435 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1519; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1521 = _fifo_in_data_T_1424 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1520; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1522 = _fifo_in_data_T_1413 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1521; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1523 = _fifo_in_data_T_1402 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1522; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1524 = _fifo_in_data_T_1391 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1523; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1525 = _fifo_in_data_T_1380 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1524; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1526 = _fifo_in_data_T_1369 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1525; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1527 = _fifo_in_data_T_1358 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1526; // @[Mux.scala 98:16]
  wire  fifo_in_valid_7 = _fifo_in_data_T_1347 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1527; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1530 = 4'h8 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1534 = _fifo_in_data_T_4 + 5'h8; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1535 = counter <= 4'h8 ? {{1'd0}, _fifo_in_data_T_1530} : _fifo_in_data_T_1534; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1537 = _fifo_in_data_T_1535 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1538 = _fifo_in_data_T_1537 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1549 = _fifo_in_data_T_1537 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1560 = _fifo_in_data_T_1537 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1571 = _fifo_in_data_T_1537 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1582 = _fifo_in_data_T_1537 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1593 = _fifo_in_data_T_1537 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1604 = _fifo_in_data_T_1537 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1615 = _fifo_in_data_T_1537 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1626 = _fifo_in_data_T_1537 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1637 = _fifo_in_data_T_1537 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1648 = _fifo_in_data_T_1537 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1659 = _fifo_in_data_T_1537 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1670 = _fifo_in_data_T_1537 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1681 = _fifo_in_data_T_1537 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1692 = _fifo_in_data_T_1537 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1703 = _fifo_in_data_T_1537 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1704 = _fifo_in_data_T_1703 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1705 = _fifo_in_data_T_1692 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1704; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1706 = _fifo_in_data_T_1681 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1705; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1707 = _fifo_in_data_T_1670 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1706; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1708 = _fifo_in_data_T_1659 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1707; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1709 = _fifo_in_data_T_1648 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1708; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1710 = _fifo_in_data_T_1637 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1709; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1711 = _fifo_in_data_T_1626 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1710; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1712 = _fifo_in_data_T_1615 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1711; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1713 = _fifo_in_data_T_1604 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1712; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1714 = _fifo_in_data_T_1593 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1713; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1715 = _fifo_in_data_T_1582 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1714; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1716 = _fifo_in_data_T_1571 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1715; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1717 = _fifo_in_data_T_1560 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1716; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1718 = _fifo_in_data_T_1549 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1717; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_8 = _fifo_in_data_T_1538 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1718; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1705 = _fifo_in_data_T_1692 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1703 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1706 = _fifo_in_data_T_1681 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1705; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1707 = _fifo_in_data_T_1670 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1706; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1708 = _fifo_in_data_T_1659 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1707; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1709 = _fifo_in_data_T_1648 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1708; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1710 = _fifo_in_data_T_1637 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1709; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1711 = _fifo_in_data_T_1626 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1710; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1712 = _fifo_in_data_T_1615 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1711; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1713 = _fifo_in_data_T_1604 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1712; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1714 = _fifo_in_data_T_1593 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1713; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1715 = _fifo_in_data_T_1582 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1714; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1716 = _fifo_in_data_T_1571 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1715; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1717 = _fifo_in_data_T_1560 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1716; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1718 = _fifo_in_data_T_1549 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1717; // @[Mux.scala 98:16]
  wire  fifo_in_valid_8 = _fifo_in_data_T_1538 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1718; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1721 = 4'h9 - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1725 = _fifo_in_data_T_4 + 5'h9; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1726 = counter <= 4'h9 ? {{1'd0}, _fifo_in_data_T_1721} : _fifo_in_data_T_1725; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1728 = _fifo_in_data_T_1726 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1729 = _fifo_in_data_T_1728 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1740 = _fifo_in_data_T_1728 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1751 = _fifo_in_data_T_1728 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1762 = _fifo_in_data_T_1728 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1773 = _fifo_in_data_T_1728 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1784 = _fifo_in_data_T_1728 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1795 = _fifo_in_data_T_1728 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1806 = _fifo_in_data_T_1728 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1817 = _fifo_in_data_T_1728 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1828 = _fifo_in_data_T_1728 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1839 = _fifo_in_data_T_1728 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1850 = _fifo_in_data_T_1728 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1861 = _fifo_in_data_T_1728 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1872 = _fifo_in_data_T_1728 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1883 = _fifo_in_data_T_1728 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1894 = _fifo_in_data_T_1728 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_1895 = _fifo_in_data_T_1894 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1896 = _fifo_in_data_T_1883 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_1895; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1897 = _fifo_in_data_T_1872 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_1896; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1898 = _fifo_in_data_T_1861 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_1897; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1899 = _fifo_in_data_T_1850 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_1898; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1900 = _fifo_in_data_T_1839 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_1899; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1901 = _fifo_in_data_T_1828 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_1900; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1902 = _fifo_in_data_T_1817 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_1901; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1903 = _fifo_in_data_T_1806 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_1902; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1904 = _fifo_in_data_T_1795 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_1903; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1905 = _fifo_in_data_T_1784 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_1904; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1906 = _fifo_in_data_T_1773 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_1905; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1907 = _fifo_in_data_T_1762 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_1906; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1908 = _fifo_in_data_T_1751 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_1907; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_1909 = _fifo_in_data_T_1740 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_1908; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_9 = _fifo_in_data_T_1729 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_1909; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1896 = _fifo_in_data_T_1883 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_1894 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1897 = _fifo_in_data_T_1872 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_1896; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1898 = _fifo_in_data_T_1861 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_1897; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1899 = _fifo_in_data_T_1850 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_1898; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1900 = _fifo_in_data_T_1839 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_1899; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1901 = _fifo_in_data_T_1828 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_1900; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1902 = _fifo_in_data_T_1817 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_1901; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1903 = _fifo_in_data_T_1806 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_1902; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1904 = _fifo_in_data_T_1795 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_1903; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1905 = _fifo_in_data_T_1784 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_1904; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1906 = _fifo_in_data_T_1773 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_1905; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1907 = _fifo_in_data_T_1762 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_1906; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1908 = _fifo_in_data_T_1751 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_1907; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_1909 = _fifo_in_data_T_1740 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_1908; // @[Mux.scala 98:16]
  wire  fifo_in_valid_9 = _fifo_in_data_T_1729 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_1909; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_1912 = 4'ha - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_1916 = _fifo_in_data_T_4 + 5'ha; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_1917 = counter <= 4'ha ? {{1'd0}, _fifo_in_data_T_1912} : _fifo_in_data_T_1916; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_1919 = _fifo_in_data_T_1917 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_1920 = _fifo_in_data_T_1919 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1931 = _fifo_in_data_T_1919 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1942 = _fifo_in_data_T_1919 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1953 = _fifo_in_data_T_1919 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1964 = _fifo_in_data_T_1919 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1975 = _fifo_in_data_T_1919 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1986 = _fifo_in_data_T_1919 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_1997 = _fifo_in_data_T_1919 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2008 = _fifo_in_data_T_1919 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2019 = _fifo_in_data_T_1919 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2030 = _fifo_in_data_T_1919 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2041 = _fifo_in_data_T_1919 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2052 = _fifo_in_data_T_1919 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2063 = _fifo_in_data_T_1919 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2074 = _fifo_in_data_T_1919 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2085 = _fifo_in_data_T_1919 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2086 = _fifo_in_data_T_2085 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2087 = _fifo_in_data_T_2074 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2086; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2088 = _fifo_in_data_T_2063 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2087; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2089 = _fifo_in_data_T_2052 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2088; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2090 = _fifo_in_data_T_2041 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2089; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2091 = _fifo_in_data_T_2030 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2090; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2092 = _fifo_in_data_T_2019 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2091; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2093 = _fifo_in_data_T_2008 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2092; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2094 = _fifo_in_data_T_1997 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2093; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2095 = _fifo_in_data_T_1986 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2094; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2096 = _fifo_in_data_T_1975 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2095; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2097 = _fifo_in_data_T_1964 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2096; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2098 = _fifo_in_data_T_1953 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2097; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2099 = _fifo_in_data_T_1942 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2098; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2100 = _fifo_in_data_T_1931 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2099; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_10 = _fifo_in_data_T_1920 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2100; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2087 = _fifo_in_data_T_2074 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2085 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2088 = _fifo_in_data_T_2063 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2087; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2089 = _fifo_in_data_T_2052 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2088; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2090 = _fifo_in_data_T_2041 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2089; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2091 = _fifo_in_data_T_2030 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2090; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2092 = _fifo_in_data_T_2019 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2091; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2093 = _fifo_in_data_T_2008 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2092; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2094 = _fifo_in_data_T_1997 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2093; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2095 = _fifo_in_data_T_1986 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2094; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2096 = _fifo_in_data_T_1975 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2095; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2097 = _fifo_in_data_T_1964 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2096; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2098 = _fifo_in_data_T_1953 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2097; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2099 = _fifo_in_data_T_1942 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2098; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2100 = _fifo_in_data_T_1931 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2099; // @[Mux.scala 98:16]
  wire  fifo_in_valid_10 = _fifo_in_data_T_1920 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2100; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2103 = 4'hb - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2107 = _fifo_in_data_T_4 + 5'hb; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_2108 = counter <= 4'hb ? {{1'd0}, _fifo_in_data_T_2103} : _fifo_in_data_T_2107; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2110 = _fifo_in_data_T_2108 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2111 = _fifo_in_data_T_2110 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2122 = _fifo_in_data_T_2110 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2133 = _fifo_in_data_T_2110 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2144 = _fifo_in_data_T_2110 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2155 = _fifo_in_data_T_2110 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2166 = _fifo_in_data_T_2110 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2177 = _fifo_in_data_T_2110 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2188 = _fifo_in_data_T_2110 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2199 = _fifo_in_data_T_2110 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2210 = _fifo_in_data_T_2110 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2221 = _fifo_in_data_T_2110 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2232 = _fifo_in_data_T_2110 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2243 = _fifo_in_data_T_2110 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2254 = _fifo_in_data_T_2110 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2265 = _fifo_in_data_T_2110 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2276 = _fifo_in_data_T_2110 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2277 = _fifo_in_data_T_2276 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2278 = _fifo_in_data_T_2265 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2277; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2279 = _fifo_in_data_T_2254 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2278; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2280 = _fifo_in_data_T_2243 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2279; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2281 = _fifo_in_data_T_2232 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2280; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2282 = _fifo_in_data_T_2221 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2281; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2283 = _fifo_in_data_T_2210 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2282; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2284 = _fifo_in_data_T_2199 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2283; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2285 = _fifo_in_data_T_2188 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2284; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2286 = _fifo_in_data_T_2177 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2285; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2287 = _fifo_in_data_T_2166 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2286; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2288 = _fifo_in_data_T_2155 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2287; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2289 = _fifo_in_data_T_2144 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2288; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2290 = _fifo_in_data_T_2133 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2289; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2291 = _fifo_in_data_T_2122 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2290; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_11 = _fifo_in_data_T_2111 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2291; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2278 = _fifo_in_data_T_2265 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2276 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2279 = _fifo_in_data_T_2254 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2278; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2280 = _fifo_in_data_T_2243 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2279; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2281 = _fifo_in_data_T_2232 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2280; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2282 = _fifo_in_data_T_2221 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2281; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2283 = _fifo_in_data_T_2210 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2282; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2284 = _fifo_in_data_T_2199 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2283; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2285 = _fifo_in_data_T_2188 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2284; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2286 = _fifo_in_data_T_2177 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2285; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2287 = _fifo_in_data_T_2166 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2286; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2288 = _fifo_in_data_T_2155 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2287; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2289 = _fifo_in_data_T_2144 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2288; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2290 = _fifo_in_data_T_2133 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2289; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2291 = _fifo_in_data_T_2122 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2290; // @[Mux.scala 98:16]
  wire  fifo_in_valid_11 = _fifo_in_data_T_2111 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2291; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2294 = 4'hc - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2298 = _fifo_in_data_T_4 + 5'hc; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_2299 = counter <= 4'hc ? {{1'd0}, _fifo_in_data_T_2294} : _fifo_in_data_T_2298; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2301 = _fifo_in_data_T_2299 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2302 = _fifo_in_data_T_2301 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2313 = _fifo_in_data_T_2301 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2324 = _fifo_in_data_T_2301 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2335 = _fifo_in_data_T_2301 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2346 = _fifo_in_data_T_2301 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2357 = _fifo_in_data_T_2301 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2368 = _fifo_in_data_T_2301 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2379 = _fifo_in_data_T_2301 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2390 = _fifo_in_data_T_2301 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2401 = _fifo_in_data_T_2301 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2412 = _fifo_in_data_T_2301 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2423 = _fifo_in_data_T_2301 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2434 = _fifo_in_data_T_2301 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2445 = _fifo_in_data_T_2301 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2456 = _fifo_in_data_T_2301 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2467 = _fifo_in_data_T_2301 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2468 = _fifo_in_data_T_2467 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2469 = _fifo_in_data_T_2456 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2468; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2470 = _fifo_in_data_T_2445 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2469; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2471 = _fifo_in_data_T_2434 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2470; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2472 = _fifo_in_data_T_2423 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2471; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2473 = _fifo_in_data_T_2412 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2472; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2474 = _fifo_in_data_T_2401 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2473; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2475 = _fifo_in_data_T_2390 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2474; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2476 = _fifo_in_data_T_2379 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2475; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2477 = _fifo_in_data_T_2368 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2476; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2478 = _fifo_in_data_T_2357 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2477; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2479 = _fifo_in_data_T_2346 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2478; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2480 = _fifo_in_data_T_2335 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2479; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2481 = _fifo_in_data_T_2324 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2480; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2482 = _fifo_in_data_T_2313 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2481; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_12 = _fifo_in_data_T_2302 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2482; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2469 = _fifo_in_data_T_2456 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2467 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2470 = _fifo_in_data_T_2445 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2469; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2471 = _fifo_in_data_T_2434 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2470; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2472 = _fifo_in_data_T_2423 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2471; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2473 = _fifo_in_data_T_2412 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2472; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2474 = _fifo_in_data_T_2401 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2473; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2475 = _fifo_in_data_T_2390 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2474; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2476 = _fifo_in_data_T_2379 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2475; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2477 = _fifo_in_data_T_2368 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2476; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2478 = _fifo_in_data_T_2357 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2477; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2479 = _fifo_in_data_T_2346 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2478; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2480 = _fifo_in_data_T_2335 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2479; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2481 = _fifo_in_data_T_2324 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2480; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2482 = _fifo_in_data_T_2313 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2481; // @[Mux.scala 98:16]
  wire  fifo_in_valid_12 = _fifo_in_data_T_2302 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2482; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2485 = 4'hd - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2489 = _fifo_in_data_T_4 + 5'hd; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_2490 = counter <= 4'hd ? {{1'd0}, _fifo_in_data_T_2485} : _fifo_in_data_T_2489; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2492 = _fifo_in_data_T_2490 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2493 = _fifo_in_data_T_2492 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2504 = _fifo_in_data_T_2492 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2515 = _fifo_in_data_T_2492 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2526 = _fifo_in_data_T_2492 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2537 = _fifo_in_data_T_2492 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2548 = _fifo_in_data_T_2492 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2559 = _fifo_in_data_T_2492 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2570 = _fifo_in_data_T_2492 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2581 = _fifo_in_data_T_2492 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2592 = _fifo_in_data_T_2492 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2603 = _fifo_in_data_T_2492 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2614 = _fifo_in_data_T_2492 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2625 = _fifo_in_data_T_2492 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2636 = _fifo_in_data_T_2492 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2647 = _fifo_in_data_T_2492 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2658 = _fifo_in_data_T_2492 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2659 = _fifo_in_data_T_2658 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2660 = _fifo_in_data_T_2647 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2659; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2661 = _fifo_in_data_T_2636 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2660; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2662 = _fifo_in_data_T_2625 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2661; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2663 = _fifo_in_data_T_2614 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2662; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2664 = _fifo_in_data_T_2603 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2663; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2665 = _fifo_in_data_T_2592 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2664; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2666 = _fifo_in_data_T_2581 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2665; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2667 = _fifo_in_data_T_2570 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2666; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2668 = _fifo_in_data_T_2559 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2667; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2669 = _fifo_in_data_T_2548 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2668; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2670 = _fifo_in_data_T_2537 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2669; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2671 = _fifo_in_data_T_2526 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2670; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2672 = _fifo_in_data_T_2515 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2671; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2673 = _fifo_in_data_T_2504 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2672; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_13 = _fifo_in_data_T_2493 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2673; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2660 = _fifo_in_data_T_2647 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2658 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2661 = _fifo_in_data_T_2636 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2660; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2662 = _fifo_in_data_T_2625 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2661; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2663 = _fifo_in_data_T_2614 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2662; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2664 = _fifo_in_data_T_2603 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2663; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2665 = _fifo_in_data_T_2592 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2664; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2666 = _fifo_in_data_T_2581 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2665; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2667 = _fifo_in_data_T_2570 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2666; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2668 = _fifo_in_data_T_2559 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2667; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2669 = _fifo_in_data_T_2548 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2668; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2670 = _fifo_in_data_T_2537 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2669; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2671 = _fifo_in_data_T_2526 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2670; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2672 = _fifo_in_data_T_2515 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2671; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2673 = _fifo_in_data_T_2504 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2672; // @[Mux.scala 98:16]
  wire  fifo_in_valid_13 = _fifo_in_data_T_2493 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2673; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2676 = 4'he - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2680 = _fifo_in_data_T_4 + 5'he; // @[BFS.scala 850:58]
  wire [4:0] _fifo_in_data_T_2681 = counter <= 4'he ? {{1'd0}, _fifo_in_data_T_2676} : _fifo_in_data_T_2680; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2683 = _fifo_in_data_T_2681 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2684 = _fifo_in_data_T_2683 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2695 = _fifo_in_data_T_2683 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2706 = _fifo_in_data_T_2683 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2717 = _fifo_in_data_T_2683 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2728 = _fifo_in_data_T_2683 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2739 = _fifo_in_data_T_2683 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2750 = _fifo_in_data_T_2683 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2761 = _fifo_in_data_T_2683 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2772 = _fifo_in_data_T_2683 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2783 = _fifo_in_data_T_2683 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2794 = _fifo_in_data_T_2683 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2805 = _fifo_in_data_T_2683 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2816 = _fifo_in_data_T_2683 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2827 = _fifo_in_data_T_2683 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2838 = _fifo_in_data_T_2683 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2849 = _fifo_in_data_T_2683 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_2850 = _fifo_in_data_T_2849 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2851 = _fifo_in_data_T_2838 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_2850; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2852 = _fifo_in_data_T_2827 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_2851; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2853 = _fifo_in_data_T_2816 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_2852; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2854 = _fifo_in_data_T_2805 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_2853; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2855 = _fifo_in_data_T_2794 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_2854; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2856 = _fifo_in_data_T_2783 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_2855; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2857 = _fifo_in_data_T_2772 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_2856; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2858 = _fifo_in_data_T_2761 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_2857; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2859 = _fifo_in_data_T_2750 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_2858; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2860 = _fifo_in_data_T_2739 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_2859; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2861 = _fifo_in_data_T_2728 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_2860; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2862 = _fifo_in_data_T_2717 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_2861; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2863 = _fifo_in_data_T_2706 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_2862; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_2864 = _fifo_in_data_T_2695 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_2863; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_14 = _fifo_in_data_T_2684 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_2864; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2851 = _fifo_in_data_T_2838 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_2849 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2852 = _fifo_in_data_T_2827 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_2851; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2853 = _fifo_in_data_T_2816 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_2852; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2854 = _fifo_in_data_T_2805 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_2853; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2855 = _fifo_in_data_T_2794 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_2854; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2856 = _fifo_in_data_T_2783 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_2855; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2857 = _fifo_in_data_T_2772 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_2856; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2858 = _fifo_in_data_T_2761 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_2857; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2859 = _fifo_in_data_T_2750 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_2858; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2860 = _fifo_in_data_T_2739 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_2859; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2861 = _fifo_in_data_T_2728 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_2860; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2862 = _fifo_in_data_T_2717 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_2861; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2863 = _fifo_in_data_T_2706 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_2862; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_2864 = _fifo_in_data_T_2695 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_2863; // @[Mux.scala 98:16]
  wire  fifo_in_valid_14 = _fifo_in_data_T_2684 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_2864; // @[Mux.scala 98:16]
  wire [3:0] _fifo_in_data_T_2867 = 4'hf - counter; // @[BFS.scala 850:34]
  wire [4:0] _fifo_in_data_T_2872 = {{1'd0}, _fifo_in_data_T_2867}; // @[BFS.scala 850:8]
  wire [4:0] _fifo_in_data_T_2874 = _fifo_in_data_T_2872 + 5'h1; // @[BFS.scala 862:39]
  wire  _fifo_in_data_T_2875 = _fifo_in_data_T_2874 == _steps_WIRE; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2886 = _fifo_in_data_T_2874 == steps_1; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2897 = _fifo_in_data_T_2874 == steps_2; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2908 = _fifo_in_data_T_2874 == steps_3; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2919 = _fifo_in_data_T_2874 == steps_4; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2930 = _fifo_in_data_T_2874 == steps_5; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2941 = _fifo_in_data_T_2874 == steps_6; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2952 = _fifo_in_data_T_2874 == steps_7; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2963 = _fifo_in_data_T_2874 == steps_8; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2974 = _fifo_in_data_T_2874 == steps_9; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2985 = _fifo_in_data_T_2874 == steps_10; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_2996 = _fifo_in_data_T_2874 == steps_11; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_3007 = _fifo_in_data_T_2874 == steps_12; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_3018 = _fifo_in_data_T_2874 == steps_13; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_3029 = _fifo_in_data_T_2874 == steps_14; // @[BFS.scala 862:46]
  wire  _fifo_in_data_T_3040 = _fifo_in_data_T_2874 == steps_15; // @[BFS.scala 862:46]
  wire [31:0] _fifo_in_data_T_3041 = _fifo_in_data_T_3040 ? in_pipeline_15_io_dout_bits_tdata : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3042 = _fifo_in_data_T_3029 ? in_pipeline_14_io_dout_bits_tdata : _fifo_in_data_T_3041; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3043 = _fifo_in_data_T_3018 ? in_pipeline_13_io_dout_bits_tdata : _fifo_in_data_T_3042; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3044 = _fifo_in_data_T_3007 ? in_pipeline_12_io_dout_bits_tdata : _fifo_in_data_T_3043; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3045 = _fifo_in_data_T_2996 ? in_pipeline_11_io_dout_bits_tdata : _fifo_in_data_T_3044; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3046 = _fifo_in_data_T_2985 ? in_pipeline_10_io_dout_bits_tdata : _fifo_in_data_T_3045; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3047 = _fifo_in_data_T_2974 ? in_pipeline_9_io_dout_bits_tdata : _fifo_in_data_T_3046; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3048 = _fifo_in_data_T_2963 ? in_pipeline_8_io_dout_bits_tdata : _fifo_in_data_T_3047; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3049 = _fifo_in_data_T_2952 ? in_pipeline_7_io_dout_bits_tdata : _fifo_in_data_T_3048; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3050 = _fifo_in_data_T_2941 ? in_pipeline_6_io_dout_bits_tdata : _fifo_in_data_T_3049; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3051 = _fifo_in_data_T_2930 ? in_pipeline_5_io_dout_bits_tdata : _fifo_in_data_T_3050; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3052 = _fifo_in_data_T_2919 ? in_pipeline_4_io_dout_bits_tdata : _fifo_in_data_T_3051; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3053 = _fifo_in_data_T_2908 ? in_pipeline_3_io_dout_bits_tdata : _fifo_in_data_T_3052; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3054 = _fifo_in_data_T_2897 ? in_pipeline_2_io_dout_bits_tdata : _fifo_in_data_T_3053; // @[Mux.scala 98:16]
  wire [31:0] _fifo_in_data_T_3055 = _fifo_in_data_T_2886 ? in_pipeline_1_io_dout_bits_tdata : _fifo_in_data_T_3054; // @[Mux.scala 98:16]
  wire [31:0] fifo_in_data_15 = _fifo_in_data_T_2875 ? in_pipeline_0_io_dout_bits_tdata : _fifo_in_data_T_3055; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3042 = _fifo_in_data_T_3029 ? in_pipeline_14_io_dout_valid : _fifo_in_data_T_3040 &
    in_pipeline_15_io_dout_valid; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3043 = _fifo_in_data_T_3018 ? in_pipeline_13_io_dout_valid : _fifo_in_valid_T_3042; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3044 = _fifo_in_data_T_3007 ? in_pipeline_12_io_dout_valid : _fifo_in_valid_T_3043; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3045 = _fifo_in_data_T_2996 ? in_pipeline_11_io_dout_valid : _fifo_in_valid_T_3044; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3046 = _fifo_in_data_T_2985 ? in_pipeline_10_io_dout_valid : _fifo_in_valid_T_3045; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3047 = _fifo_in_data_T_2974 ? in_pipeline_9_io_dout_valid : _fifo_in_valid_T_3046; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3048 = _fifo_in_data_T_2963 ? in_pipeline_8_io_dout_valid : _fifo_in_valid_T_3047; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3049 = _fifo_in_data_T_2952 ? in_pipeline_7_io_dout_valid : _fifo_in_valid_T_3048; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3050 = _fifo_in_data_T_2941 ? in_pipeline_6_io_dout_valid : _fifo_in_valid_T_3049; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3051 = _fifo_in_data_T_2930 ? in_pipeline_5_io_dout_valid : _fifo_in_valid_T_3050; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3052 = _fifo_in_data_T_2919 ? in_pipeline_4_io_dout_valid : _fifo_in_valid_T_3051; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3053 = _fifo_in_data_T_2908 ? in_pipeline_3_io_dout_valid : _fifo_in_valid_T_3052; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3054 = _fifo_in_data_T_2897 ? in_pipeline_2_io_dout_valid : _fifo_in_valid_T_3053; // @[Mux.scala 98:16]
  wire  _fifo_in_valid_T_3055 = _fifo_in_data_T_2886 ? in_pipeline_1_io_dout_valid : _fifo_in_valid_T_3054; // @[Mux.scala 98:16]
  wire  fifo_in_valid_15 = _fifo_in_data_T_2875 ? in_pipeline_0_io_dout_valid : _fifo_in_valid_T_3055; // @[Mux.scala 98:16]
  wire [31:0] collector_data_1 = collector_fifos_1_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_0 = collector_fifos_0_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_3 = collector_fifos_3_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_2 = collector_fifos_2_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_5 = collector_fifos_5_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_4 = collector_fifos_4_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_7 = collector_fifos_7_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_6 = collector_fifos_6_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [255:0] io_out_dout_lo = {collector_data_7,collector_data_6,collector_data_5,collector_data_4,collector_data_3,
    collector_data_2,collector_data_1,collector_data_0}; // @[BFS.scala 877:39]
  wire [31:0] collector_data_9 = collector_fifos_9_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_8 = collector_fifos_8_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_11 = collector_fifos_11_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_10 = collector_fifos_10_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_13 = collector_fifos_13_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_12 = collector_fifos_12_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_15 = collector_fifos_15_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [31:0] collector_data_14 = collector_fifos_14_dout; // @[BFS.scala 830:28 BFS.scala 869:25]
  wire [255:0] io_out_dout_hi = {collector_data_15,collector_data_14,collector_data_13,collector_data_12,
    collector_data_11,collector_data_10,collector_data_9,collector_data_8}; // @[BFS.scala 877:39]
  wire [8:0] _io_out_data_count_WIRE = {{4'd0}, collector_fifos_0_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_WIRE_1 = {{4'd0}, collector_fifos_1_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_1 = _io_out_data_count_WIRE + _io_out_data_count_WIRE_1; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_2 = {{4'd0}, collector_fifos_2_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_3 = _io_out_data_count_T_1 + _io_out_data_count_WIRE_2; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_3 = {{4'd0}, collector_fifos_3_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_5 = _io_out_data_count_T_3 + _io_out_data_count_WIRE_3; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_4 = {{4'd0}, collector_fifos_4_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_7 = _io_out_data_count_T_5 + _io_out_data_count_WIRE_4; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_5 = {{4'd0}, collector_fifos_5_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_9 = _io_out_data_count_T_7 + _io_out_data_count_WIRE_5; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_6 = {{4'd0}, collector_fifos_6_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_11 = _io_out_data_count_T_9 + _io_out_data_count_WIRE_6; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_7 = {{4'd0}, collector_fifos_7_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_13 = _io_out_data_count_T_11 + _io_out_data_count_WIRE_7; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_8 = {{4'd0}, collector_fifos_8_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_15 = _io_out_data_count_T_13 + _io_out_data_count_WIRE_8; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_9 = {{4'd0}, collector_fifos_9_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_17 = _io_out_data_count_T_15 + _io_out_data_count_WIRE_9; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_10 = {{4'd0}, collector_fifos_10_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_19 = _io_out_data_count_T_17 + _io_out_data_count_WIRE_10; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_11 = {{4'd0}, collector_fifos_11_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_21 = _io_out_data_count_T_19 + _io_out_data_count_WIRE_11; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_12 = {{4'd0}, collector_fifos_12_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_23 = _io_out_data_count_T_21 + _io_out_data_count_WIRE_12; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_13 = {{4'd0}, collector_fifos_13_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_25 = _io_out_data_count_T_23 + _io_out_data_count_WIRE_13; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_14 = {{4'd0}, collector_fifos_14_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  wire [8:0] _io_out_data_count_T_27 = _io_out_data_count_T_25 + _io_out_data_count_WIRE_14; // @[BFS.scala 878:134]
  wire [8:0] _io_out_data_count_WIRE_15 = {{4'd0}, collector_fifos_15_data_count}; // @[BFS.scala 878:73 BFS.scala 878:73]
  collector_fifo_0 collector_fifos_0 ( // @[BFS.scala 826:16]
    .full(collector_fifos_0_full),
    .din(collector_fifos_0_din),
    .wr_en(collector_fifos_0_wr_en),
    .empty(collector_fifos_0_empty),
    .dout(collector_fifos_0_dout),
    .rd_en(collector_fifos_0_rd_en),
    .data_count(collector_fifos_0_data_count),
    .clk(collector_fifos_0_clk),
    .srst(collector_fifos_0_srst),
    .valid(collector_fifos_0_valid)
  );
  collector_fifo_0 collector_fifos_1 ( // @[BFS.scala 826:16]
    .full(collector_fifos_1_full),
    .din(collector_fifos_1_din),
    .wr_en(collector_fifos_1_wr_en),
    .empty(collector_fifos_1_empty),
    .dout(collector_fifos_1_dout),
    .rd_en(collector_fifos_1_rd_en),
    .data_count(collector_fifos_1_data_count),
    .clk(collector_fifos_1_clk),
    .srst(collector_fifos_1_srst),
    .valid(collector_fifos_1_valid)
  );
  collector_fifo_0 collector_fifos_2 ( // @[BFS.scala 826:16]
    .full(collector_fifos_2_full),
    .din(collector_fifos_2_din),
    .wr_en(collector_fifos_2_wr_en),
    .empty(collector_fifos_2_empty),
    .dout(collector_fifos_2_dout),
    .rd_en(collector_fifos_2_rd_en),
    .data_count(collector_fifos_2_data_count),
    .clk(collector_fifos_2_clk),
    .srst(collector_fifos_2_srst),
    .valid(collector_fifos_2_valid)
  );
  collector_fifo_0 collector_fifos_3 ( // @[BFS.scala 826:16]
    .full(collector_fifos_3_full),
    .din(collector_fifos_3_din),
    .wr_en(collector_fifos_3_wr_en),
    .empty(collector_fifos_3_empty),
    .dout(collector_fifos_3_dout),
    .rd_en(collector_fifos_3_rd_en),
    .data_count(collector_fifos_3_data_count),
    .clk(collector_fifos_3_clk),
    .srst(collector_fifos_3_srst),
    .valid(collector_fifos_3_valid)
  );
  collector_fifo_0 collector_fifos_4 ( // @[BFS.scala 826:16]
    .full(collector_fifos_4_full),
    .din(collector_fifos_4_din),
    .wr_en(collector_fifos_4_wr_en),
    .empty(collector_fifos_4_empty),
    .dout(collector_fifos_4_dout),
    .rd_en(collector_fifos_4_rd_en),
    .data_count(collector_fifos_4_data_count),
    .clk(collector_fifos_4_clk),
    .srst(collector_fifos_4_srst),
    .valid(collector_fifos_4_valid)
  );
  collector_fifo_0 collector_fifos_5 ( // @[BFS.scala 826:16]
    .full(collector_fifos_5_full),
    .din(collector_fifos_5_din),
    .wr_en(collector_fifos_5_wr_en),
    .empty(collector_fifos_5_empty),
    .dout(collector_fifos_5_dout),
    .rd_en(collector_fifos_5_rd_en),
    .data_count(collector_fifos_5_data_count),
    .clk(collector_fifos_5_clk),
    .srst(collector_fifos_5_srst),
    .valid(collector_fifos_5_valid)
  );
  collector_fifo_0 collector_fifos_6 ( // @[BFS.scala 826:16]
    .full(collector_fifos_6_full),
    .din(collector_fifos_6_din),
    .wr_en(collector_fifos_6_wr_en),
    .empty(collector_fifos_6_empty),
    .dout(collector_fifos_6_dout),
    .rd_en(collector_fifos_6_rd_en),
    .data_count(collector_fifos_6_data_count),
    .clk(collector_fifos_6_clk),
    .srst(collector_fifos_6_srst),
    .valid(collector_fifos_6_valid)
  );
  collector_fifo_0 collector_fifos_7 ( // @[BFS.scala 826:16]
    .full(collector_fifos_7_full),
    .din(collector_fifos_7_din),
    .wr_en(collector_fifos_7_wr_en),
    .empty(collector_fifos_7_empty),
    .dout(collector_fifos_7_dout),
    .rd_en(collector_fifos_7_rd_en),
    .data_count(collector_fifos_7_data_count),
    .clk(collector_fifos_7_clk),
    .srst(collector_fifos_7_srst),
    .valid(collector_fifos_7_valid)
  );
  collector_fifo_0 collector_fifos_8 ( // @[BFS.scala 826:16]
    .full(collector_fifos_8_full),
    .din(collector_fifos_8_din),
    .wr_en(collector_fifos_8_wr_en),
    .empty(collector_fifos_8_empty),
    .dout(collector_fifos_8_dout),
    .rd_en(collector_fifos_8_rd_en),
    .data_count(collector_fifos_8_data_count),
    .clk(collector_fifos_8_clk),
    .srst(collector_fifos_8_srst),
    .valid(collector_fifos_8_valid)
  );
  collector_fifo_0 collector_fifos_9 ( // @[BFS.scala 826:16]
    .full(collector_fifos_9_full),
    .din(collector_fifos_9_din),
    .wr_en(collector_fifos_9_wr_en),
    .empty(collector_fifos_9_empty),
    .dout(collector_fifos_9_dout),
    .rd_en(collector_fifos_9_rd_en),
    .data_count(collector_fifos_9_data_count),
    .clk(collector_fifos_9_clk),
    .srst(collector_fifos_9_srst),
    .valid(collector_fifos_9_valid)
  );
  collector_fifo_0 collector_fifos_10 ( // @[BFS.scala 826:16]
    .full(collector_fifos_10_full),
    .din(collector_fifos_10_din),
    .wr_en(collector_fifos_10_wr_en),
    .empty(collector_fifos_10_empty),
    .dout(collector_fifos_10_dout),
    .rd_en(collector_fifos_10_rd_en),
    .data_count(collector_fifos_10_data_count),
    .clk(collector_fifos_10_clk),
    .srst(collector_fifos_10_srst),
    .valid(collector_fifos_10_valid)
  );
  collector_fifo_0 collector_fifos_11 ( // @[BFS.scala 826:16]
    .full(collector_fifos_11_full),
    .din(collector_fifos_11_din),
    .wr_en(collector_fifos_11_wr_en),
    .empty(collector_fifos_11_empty),
    .dout(collector_fifos_11_dout),
    .rd_en(collector_fifos_11_rd_en),
    .data_count(collector_fifos_11_data_count),
    .clk(collector_fifos_11_clk),
    .srst(collector_fifos_11_srst),
    .valid(collector_fifos_11_valid)
  );
  collector_fifo_0 collector_fifos_12 ( // @[BFS.scala 826:16]
    .full(collector_fifos_12_full),
    .din(collector_fifos_12_din),
    .wr_en(collector_fifos_12_wr_en),
    .empty(collector_fifos_12_empty),
    .dout(collector_fifos_12_dout),
    .rd_en(collector_fifos_12_rd_en),
    .data_count(collector_fifos_12_data_count),
    .clk(collector_fifos_12_clk),
    .srst(collector_fifos_12_srst),
    .valid(collector_fifos_12_valid)
  );
  collector_fifo_0 collector_fifos_13 ( // @[BFS.scala 826:16]
    .full(collector_fifos_13_full),
    .din(collector_fifos_13_din),
    .wr_en(collector_fifos_13_wr_en),
    .empty(collector_fifos_13_empty),
    .dout(collector_fifos_13_dout),
    .rd_en(collector_fifos_13_rd_en),
    .data_count(collector_fifos_13_data_count),
    .clk(collector_fifos_13_clk),
    .srst(collector_fifos_13_srst),
    .valid(collector_fifos_13_valid)
  );
  collector_fifo_0 collector_fifos_14 ( // @[BFS.scala 826:16]
    .full(collector_fifos_14_full),
    .din(collector_fifos_14_din),
    .wr_en(collector_fifos_14_wr_en),
    .empty(collector_fifos_14_empty),
    .dout(collector_fifos_14_dout),
    .rd_en(collector_fifos_14_rd_en),
    .data_count(collector_fifos_14_data_count),
    .clk(collector_fifos_14_clk),
    .srst(collector_fifos_14_srst),
    .valid(collector_fifos_14_valid)
  );
  collector_fifo_0 collector_fifos_15 ( // @[BFS.scala 826:16]
    .full(collector_fifos_15_full),
    .din(collector_fifos_15_din),
    .wr_en(collector_fifos_15_wr_en),
    .empty(collector_fifos_15_empty),
    .dout(collector_fifos_15_dout),
    .rd_en(collector_fifos_15_rd_en),
    .data_count(collector_fifos_15_data_count),
    .clk(collector_fifos_15_clk),
    .srst(collector_fifos_15_srst),
    .valid(collector_fifos_15_valid)
  );
  pipeline in_pipeline_0 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_0_clock),
    .reset(in_pipeline_0_reset),
    .io_dout_ready(in_pipeline_0_io_dout_ready),
    .io_dout_valid(in_pipeline_0_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_0_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_0_io_din_ready),
    .io_din_valid(in_pipeline_0_io_din_valid),
    .io_din_bits_tdata(in_pipeline_0_io_din_bits_tdata)
  );
  pipeline in_pipeline_1 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_1_clock),
    .reset(in_pipeline_1_reset),
    .io_dout_ready(in_pipeline_1_io_dout_ready),
    .io_dout_valid(in_pipeline_1_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_1_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_1_io_din_ready),
    .io_din_valid(in_pipeline_1_io_din_valid),
    .io_din_bits_tdata(in_pipeline_1_io_din_bits_tdata)
  );
  pipeline in_pipeline_2 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_2_clock),
    .reset(in_pipeline_2_reset),
    .io_dout_ready(in_pipeline_2_io_dout_ready),
    .io_dout_valid(in_pipeline_2_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_2_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_2_io_din_ready),
    .io_din_valid(in_pipeline_2_io_din_valid),
    .io_din_bits_tdata(in_pipeline_2_io_din_bits_tdata)
  );
  pipeline in_pipeline_3 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_3_clock),
    .reset(in_pipeline_3_reset),
    .io_dout_ready(in_pipeline_3_io_dout_ready),
    .io_dout_valid(in_pipeline_3_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_3_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_3_io_din_ready),
    .io_din_valid(in_pipeline_3_io_din_valid),
    .io_din_bits_tdata(in_pipeline_3_io_din_bits_tdata)
  );
  pipeline in_pipeline_4 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_4_clock),
    .reset(in_pipeline_4_reset),
    .io_dout_ready(in_pipeline_4_io_dout_ready),
    .io_dout_valid(in_pipeline_4_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_4_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_4_io_din_ready),
    .io_din_valid(in_pipeline_4_io_din_valid),
    .io_din_bits_tdata(in_pipeline_4_io_din_bits_tdata)
  );
  pipeline in_pipeline_5 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_5_clock),
    .reset(in_pipeline_5_reset),
    .io_dout_ready(in_pipeline_5_io_dout_ready),
    .io_dout_valid(in_pipeline_5_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_5_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_5_io_din_ready),
    .io_din_valid(in_pipeline_5_io_din_valid),
    .io_din_bits_tdata(in_pipeline_5_io_din_bits_tdata)
  );
  pipeline in_pipeline_6 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_6_clock),
    .reset(in_pipeline_6_reset),
    .io_dout_ready(in_pipeline_6_io_dout_ready),
    .io_dout_valid(in_pipeline_6_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_6_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_6_io_din_ready),
    .io_din_valid(in_pipeline_6_io_din_valid),
    .io_din_bits_tdata(in_pipeline_6_io_din_bits_tdata)
  );
  pipeline in_pipeline_7 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_7_clock),
    .reset(in_pipeline_7_reset),
    .io_dout_ready(in_pipeline_7_io_dout_ready),
    .io_dout_valid(in_pipeline_7_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_7_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_7_io_din_ready),
    .io_din_valid(in_pipeline_7_io_din_valid),
    .io_din_bits_tdata(in_pipeline_7_io_din_bits_tdata)
  );
  pipeline in_pipeline_8 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_8_clock),
    .reset(in_pipeline_8_reset),
    .io_dout_ready(in_pipeline_8_io_dout_ready),
    .io_dout_valid(in_pipeline_8_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_8_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_8_io_din_ready),
    .io_din_valid(in_pipeline_8_io_din_valid),
    .io_din_bits_tdata(in_pipeline_8_io_din_bits_tdata)
  );
  pipeline in_pipeline_9 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_9_clock),
    .reset(in_pipeline_9_reset),
    .io_dout_ready(in_pipeline_9_io_dout_ready),
    .io_dout_valid(in_pipeline_9_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_9_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_9_io_din_ready),
    .io_din_valid(in_pipeline_9_io_din_valid),
    .io_din_bits_tdata(in_pipeline_9_io_din_bits_tdata)
  );
  pipeline in_pipeline_10 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_10_clock),
    .reset(in_pipeline_10_reset),
    .io_dout_ready(in_pipeline_10_io_dout_ready),
    .io_dout_valid(in_pipeline_10_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_10_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_10_io_din_ready),
    .io_din_valid(in_pipeline_10_io_din_valid),
    .io_din_bits_tdata(in_pipeline_10_io_din_bits_tdata)
  );
  pipeline in_pipeline_11 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_11_clock),
    .reset(in_pipeline_11_reset),
    .io_dout_ready(in_pipeline_11_io_dout_ready),
    .io_dout_valid(in_pipeline_11_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_11_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_11_io_din_ready),
    .io_din_valid(in_pipeline_11_io_din_valid),
    .io_din_bits_tdata(in_pipeline_11_io_din_bits_tdata)
  );
  pipeline in_pipeline_12 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_12_clock),
    .reset(in_pipeline_12_reset),
    .io_dout_ready(in_pipeline_12_io_dout_ready),
    .io_dout_valid(in_pipeline_12_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_12_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_12_io_din_ready),
    .io_din_valid(in_pipeline_12_io_din_valid),
    .io_din_bits_tdata(in_pipeline_12_io_din_bits_tdata)
  );
  pipeline in_pipeline_13 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_13_clock),
    .reset(in_pipeline_13_reset),
    .io_dout_ready(in_pipeline_13_io_dout_ready),
    .io_dout_valid(in_pipeline_13_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_13_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_13_io_din_ready),
    .io_din_valid(in_pipeline_13_io_din_valid),
    .io_din_bits_tdata(in_pipeline_13_io_din_bits_tdata)
  );
  pipeline in_pipeline_14 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_14_clock),
    .reset(in_pipeline_14_reset),
    .io_dout_ready(in_pipeline_14_io_dout_ready),
    .io_dout_valid(in_pipeline_14_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_14_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_14_io_din_ready),
    .io_din_valid(in_pipeline_14_io_din_valid),
    .io_din_bits_tdata(in_pipeline_14_io_din_bits_tdata)
  );
  pipeline in_pipeline_15 ( // @[BFS.scala 832:11]
    .clock(in_pipeline_15_clock),
    .reset(in_pipeline_15_reset),
    .io_dout_ready(in_pipeline_15_io_dout_ready),
    .io_dout_valid(in_pipeline_15_io_dout_valid),
    .io_dout_bits_tdata(in_pipeline_15_io_dout_bits_tdata),
    .io_din_ready(in_pipeline_15_io_din_ready),
    .io_din_valid(in_pipeline_15_io_din_valid),
    .io_din_bits_tdata(in_pipeline_15_io_din_bits_tdata)
  );
  assign io_in_0_ready = in_pipeline_0_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_1_ready = in_pipeline_1_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_2_ready = in_pipeline_2_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_3_ready = in_pipeline_3_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_4_ready = in_pipeline_4_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_5_ready = in_pipeline_5_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_6_ready = in_pipeline_6_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_7_ready = in_pipeline_7_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_8_ready = in_pipeline_8_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_9_ready = in_pipeline_9_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_10_ready = in_pipeline_10_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_11_ready = in_pipeline_11_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_12_ready = in_pipeline_12_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_13_ready = in_pipeline_13_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_14_ready = in_pipeline_14_io_din_ready; // @[BFS.scala 836:16]
  assign io_in_15_ready = in_pipeline_15_io_din_ready; // @[BFS.scala 836:16]
  assign io_out_full = ~fifos_ready; // @[BFS.scala 879:18]
  assign io_out_dout = {io_out_dout_hi,io_out_dout_lo}; // @[BFS.scala 877:39]
  assign io_out_data_count = _io_out_data_count_T_27 + _io_out_data_count_WIRE_15; // @[BFS.scala 878:134]
  assign io_out_valid = collector_fifos_0_valid | collector_fifos_1_valid | collector_fifos_2_valid |
    collector_fifos_3_valid | collector_fifos_4_valid | collector_fifos_5_valid | collector_fifos_6_valid |
    collector_fifos_7_valid | collector_fifos_8_valid | collector_fifos_9_valid | collector_fifos_10_valid |
    collector_fifos_11_valid | collector_fifos_12_valid | collector_fifos_13_valid | collector_fifos_14_valid |
    collector_fifos_15_valid; // @[BFS.scala 876:80]
  assign collector_fifos_0_din = io_is_current_tier ? io_out_din[31:0] : fifo_in_data; // @[BFS.scala 867:22]
  assign collector_fifos_0_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid; // @[BFS.scala 868:24]
  assign collector_fifos_0_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_0_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_0_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_1_din = io_is_current_tier ? io_out_din[63:32] : fifo_in_data_1; // @[BFS.scala 867:22]
  assign collector_fifos_1_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_1; // @[BFS.scala 868:24]
  assign collector_fifos_1_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_1_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_1_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_2_din = io_is_current_tier ? io_out_din[95:64] : fifo_in_data_2; // @[BFS.scala 867:22]
  assign collector_fifos_2_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_2; // @[BFS.scala 868:24]
  assign collector_fifos_2_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_2_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_2_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_3_din = io_is_current_tier ? io_out_din[127:96] : fifo_in_data_3; // @[BFS.scala 867:22]
  assign collector_fifos_3_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_3; // @[BFS.scala 868:24]
  assign collector_fifos_3_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_3_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_3_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_4_din = io_is_current_tier ? io_out_din[159:128] : fifo_in_data_4; // @[BFS.scala 867:22]
  assign collector_fifos_4_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_4; // @[BFS.scala 868:24]
  assign collector_fifos_4_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_4_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_4_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_5_din = io_is_current_tier ? io_out_din[191:160] : fifo_in_data_5; // @[BFS.scala 867:22]
  assign collector_fifos_5_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_5; // @[BFS.scala 868:24]
  assign collector_fifos_5_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_5_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_5_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_6_din = io_is_current_tier ? io_out_din[223:192] : fifo_in_data_6; // @[BFS.scala 867:22]
  assign collector_fifos_6_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_6; // @[BFS.scala 868:24]
  assign collector_fifos_6_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_6_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_6_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_7_din = io_is_current_tier ? io_out_din[255:224] : fifo_in_data_7; // @[BFS.scala 867:22]
  assign collector_fifos_7_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_7; // @[BFS.scala 868:24]
  assign collector_fifos_7_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_7_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_7_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_8_din = io_is_current_tier ? io_out_din[287:256] : fifo_in_data_8; // @[BFS.scala 867:22]
  assign collector_fifos_8_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_8; // @[BFS.scala 868:24]
  assign collector_fifos_8_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_8_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_8_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_9_din = io_is_current_tier ? io_out_din[319:288] : fifo_in_data_9; // @[BFS.scala 867:22]
  assign collector_fifos_9_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_9; // @[BFS.scala 868:24]
  assign collector_fifos_9_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_9_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_9_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_10_din = io_is_current_tier ? io_out_din[351:320] : fifo_in_data_10; // @[BFS.scala 867:22]
  assign collector_fifos_10_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_10; // @[BFS.scala 868:24]
  assign collector_fifos_10_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_10_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_10_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_11_din = io_is_current_tier ? io_out_din[383:352] : fifo_in_data_11; // @[BFS.scala 867:22]
  assign collector_fifos_11_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_11; // @[BFS.scala 868:24]
  assign collector_fifos_11_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_11_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_11_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_12_din = io_is_current_tier ? io_out_din[415:384] : fifo_in_data_12; // @[BFS.scala 867:22]
  assign collector_fifos_12_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_12; // @[BFS.scala 868:24]
  assign collector_fifos_12_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_12_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_12_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_13_din = io_is_current_tier ? io_out_din[447:416] : fifo_in_data_13; // @[BFS.scala 867:22]
  assign collector_fifos_13_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_13; // @[BFS.scala 868:24]
  assign collector_fifos_13_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_13_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_13_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_14_din = io_is_current_tier ? io_out_din[479:448] : fifo_in_data_14; // @[BFS.scala 867:22]
  assign collector_fifos_14_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_14; // @[BFS.scala 868:24]
  assign collector_fifos_14_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_14_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_14_srst = reset; // @[BFS.scala 871:32]
  assign collector_fifos_15_din = io_is_current_tier ? io_out_din[511:480] : fifo_in_data_15; // @[BFS.scala 867:22]
  assign collector_fifos_15_wr_en = io_is_current_tier ? io_out_wr_en : fifo_in_valid_15; // @[BFS.scala 868:24]
  assign collector_fifos_15_rd_en = io_out_rd_en; // @[BFS.scala 872:18]
  assign collector_fifos_15_clk = clock; // @[BFS.scala 870:31]
  assign collector_fifos_15_srst = reset; // @[BFS.scala 871:32]
  assign in_pipeline_0_clock = clock;
  assign in_pipeline_0_reset = reset;
  assign in_pipeline_0_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_0_io_din_valid = io_in_0_valid; // @[BFS.scala 836:16]
  assign in_pipeline_0_io_din_bits_tdata = io_in_0_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_1_clock = clock;
  assign in_pipeline_1_reset = reset;
  assign in_pipeline_1_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_1_io_din_valid = io_in_1_valid; // @[BFS.scala 836:16]
  assign in_pipeline_1_io_din_bits_tdata = io_in_1_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_2_clock = clock;
  assign in_pipeline_2_reset = reset;
  assign in_pipeline_2_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_2_io_din_valid = io_in_2_valid; // @[BFS.scala 836:16]
  assign in_pipeline_2_io_din_bits_tdata = io_in_2_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_3_clock = clock;
  assign in_pipeline_3_reset = reset;
  assign in_pipeline_3_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_3_io_din_valid = io_in_3_valid; // @[BFS.scala 836:16]
  assign in_pipeline_3_io_din_bits_tdata = io_in_3_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_4_clock = clock;
  assign in_pipeline_4_reset = reset;
  assign in_pipeline_4_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_4_io_din_valid = io_in_4_valid; // @[BFS.scala 836:16]
  assign in_pipeline_4_io_din_bits_tdata = io_in_4_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_5_clock = clock;
  assign in_pipeline_5_reset = reset;
  assign in_pipeline_5_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_5_io_din_valid = io_in_5_valid; // @[BFS.scala 836:16]
  assign in_pipeline_5_io_din_bits_tdata = io_in_5_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_6_clock = clock;
  assign in_pipeline_6_reset = reset;
  assign in_pipeline_6_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_6_io_din_valid = io_in_6_valid; // @[BFS.scala 836:16]
  assign in_pipeline_6_io_din_bits_tdata = io_in_6_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_7_clock = clock;
  assign in_pipeline_7_reset = reset;
  assign in_pipeline_7_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_7_io_din_valid = io_in_7_valid; // @[BFS.scala 836:16]
  assign in_pipeline_7_io_din_bits_tdata = io_in_7_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_8_clock = clock;
  assign in_pipeline_8_reset = reset;
  assign in_pipeline_8_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_8_io_din_valid = io_in_8_valid; // @[BFS.scala 836:16]
  assign in_pipeline_8_io_din_bits_tdata = io_in_8_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_9_clock = clock;
  assign in_pipeline_9_reset = reset;
  assign in_pipeline_9_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_9_io_din_valid = io_in_9_valid; // @[BFS.scala 836:16]
  assign in_pipeline_9_io_din_bits_tdata = io_in_9_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_10_clock = clock;
  assign in_pipeline_10_reset = reset;
  assign in_pipeline_10_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_10_io_din_valid = io_in_10_valid; // @[BFS.scala 836:16]
  assign in_pipeline_10_io_din_bits_tdata = io_in_10_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_11_clock = clock;
  assign in_pipeline_11_reset = reset;
  assign in_pipeline_11_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_11_io_din_valid = io_in_11_valid; // @[BFS.scala 836:16]
  assign in_pipeline_11_io_din_bits_tdata = io_in_11_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_12_clock = clock;
  assign in_pipeline_12_reset = reset;
  assign in_pipeline_12_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_12_io_din_valid = io_in_12_valid; // @[BFS.scala 836:16]
  assign in_pipeline_12_io_din_bits_tdata = io_in_12_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_13_clock = clock;
  assign in_pipeline_13_reset = reset;
  assign in_pipeline_13_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_13_io_din_valid = io_in_13_valid; // @[BFS.scala 836:16]
  assign in_pipeline_13_io_din_bits_tdata = io_in_13_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_14_clock = clock;
  assign in_pipeline_14_reset = reset;
  assign in_pipeline_14_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_14_io_din_valid = io_in_14_valid; // @[BFS.scala 836:16]
  assign in_pipeline_14_io_din_bits_tdata = io_in_14_bits_tdata; // @[BFS.scala 836:16]
  assign in_pipeline_15_clock = clock;
  assign in_pipeline_15_reset = reset;
  assign in_pipeline_15_io_dout_ready = io_is_current_tier ? 1'h0 : fifos_ready; // @[BFS.scala 837:29]
  assign in_pipeline_15_io_din_valid = io_in_15_valid; // @[BFS.scala 836:16]
  assign in_pipeline_15_io_din_bits_tdata = io_in_15_bits_tdata; // @[BFS.scala 836:16]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 829:24]
      counter <= 4'h0; // @[BFS.scala 829:24]
    end else begin
      counter <= _GEN_1[3:0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multi_port_mc(
  input          clock,
  input          reset,
  input          io_cacheable_out_ready,
  output         io_cacheable_out_valid,
  output [511:0] io_cacheable_out_bits_tdata,
  output [15:0]  io_cacheable_out_bits_tkeep,
  output         io_cacheable_in_0_ready,
  input          io_cacheable_in_0_valid,
  input  [31:0]  io_cacheable_in_0_bits_tdata,
  output         io_cacheable_in_1_ready,
  input          io_cacheable_in_1_valid,
  input  [31:0]  io_cacheable_in_1_bits_tdata,
  output         io_cacheable_in_2_ready,
  input          io_cacheable_in_2_valid,
  input  [31:0]  io_cacheable_in_2_bits_tdata,
  output         io_cacheable_in_3_ready,
  input          io_cacheable_in_3_valid,
  input  [31:0]  io_cacheable_in_3_bits_tdata,
  output         io_cacheable_in_4_ready,
  input          io_cacheable_in_4_valid,
  input  [31:0]  io_cacheable_in_4_bits_tdata,
  output         io_cacheable_in_5_ready,
  input          io_cacheable_in_5_valid,
  input  [31:0]  io_cacheable_in_5_bits_tdata,
  output         io_cacheable_in_6_ready,
  input          io_cacheable_in_6_valid,
  input  [31:0]  io_cacheable_in_6_bits_tdata,
  output         io_cacheable_in_7_ready,
  input          io_cacheable_in_7_valid,
  input  [31:0]  io_cacheable_in_7_bits_tdata,
  output         io_cacheable_in_8_ready,
  input          io_cacheable_in_8_valid,
  input  [31:0]  io_cacheable_in_8_bits_tdata,
  output         io_cacheable_in_9_ready,
  input          io_cacheable_in_9_valid,
  input  [31:0]  io_cacheable_in_9_bits_tdata,
  output         io_cacheable_in_10_ready,
  input          io_cacheable_in_10_valid,
  input  [31:0]  io_cacheable_in_10_bits_tdata,
  output         io_cacheable_in_11_ready,
  input          io_cacheable_in_11_valid,
  input  [31:0]  io_cacheable_in_11_bits_tdata,
  output         io_cacheable_in_12_ready,
  input          io_cacheable_in_12_valid,
  input  [31:0]  io_cacheable_in_12_bits_tdata,
  output         io_cacheable_in_13_ready,
  input          io_cacheable_in_13_valid,
  input  [31:0]  io_cacheable_in_13_bits_tdata,
  output         io_cacheable_in_14_ready,
  input          io_cacheable_in_14_valid,
  input  [31:0]  io_cacheable_in_14_bits_tdata,
  output         io_cacheable_in_15_ready,
  input          io_cacheable_in_15_valid,
  input  [31:0]  io_cacheable_in_15_bits_tdata,
  output         io_non_cacheable_in_aw_ready,
  input          io_non_cacheable_in_aw_valid,
  input  [63:0]  io_non_cacheable_in_aw_bits_awaddr,
  input  [6:0]   io_non_cacheable_in_aw_bits_awid,
  output         io_non_cacheable_in_w_ready,
  input          io_non_cacheable_in_w_valid,
  input  [511:0] io_non_cacheable_in_w_bits_wdata,
  input  [63:0]  io_non_cacheable_in_w_bits_wstrb,
  input          io_ddr_out_0_aw_ready,
  output         io_ddr_out_0_aw_valid,
  output [63:0]  io_ddr_out_0_aw_bits_awaddr,
  input          io_ddr_out_0_ar_ready,
  output         io_ddr_out_0_ar_valid,
  output [63:0]  io_ddr_out_0_ar_bits_araddr,
  input          io_ddr_out_0_w_ready,
  output         io_ddr_out_0_w_valid,
  output [511:0] io_ddr_out_0_w_bits_wdata,
  output         io_ddr_out_0_w_bits_wlast,
  input          io_ddr_out_0_r_valid,
  input  [511:0] io_ddr_out_0_r_bits_rdata,
  input          io_ddr_out_0_r_bits_rlast,
  input          io_ddr_out_1_aw_ready,
  output         io_ddr_out_1_aw_valid,
  output [63:0]  io_ddr_out_1_aw_bits_awaddr,
  output [6:0]   io_ddr_out_1_aw_bits_awid,
  input          io_ddr_out_1_w_ready,
  output         io_ddr_out_1_w_valid,
  output [511:0] io_ddr_out_1_w_bits_wdata,
  output [63:0]  io_ddr_out_1_w_bits_wstrb,
  input  [63:0]  io_tiers_base_addr_0,
  input  [63:0]  io_tiers_base_addr_1,
  output [31:0]  io_unvisited_size,
  input          io_start,
  input          io_signal,
  input          io_end,
  output         io_signal_ack
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  tier_fifo_0_clock; // @[BFS.scala 903:46]
  wire  tier_fifo_0_reset; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_0_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_0_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_0_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_1_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_1_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_1_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_2_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_2_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_2_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_3_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_3_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_3_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_4_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_4_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_4_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_5_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_5_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_5_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_6_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_6_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_6_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_7_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_7_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_7_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_8_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_8_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_8_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_9_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_9_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_9_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_10_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_10_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_10_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_11_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_11_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_11_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_12_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_12_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_12_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_13_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_13_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_13_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_14_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_14_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_14_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_15_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_in_15_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_0_io_in_15_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_out_full; // @[BFS.scala 903:46]
  wire [511:0] tier_fifo_0_io_out_din; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_out_wr_en; // @[BFS.scala 903:46]
  wire [511:0] tier_fifo_0_io_out_dout; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_out_rd_en; // @[BFS.scala 903:46]
  wire [8:0] tier_fifo_0_io_out_data_count; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_out_valid; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_flush; // @[BFS.scala 903:46]
  wire  tier_fifo_0_io_is_current_tier; // @[BFS.scala 903:46]
  wire  tier_fifo_1_clock; // @[BFS.scala 903:46]
  wire  tier_fifo_1_reset; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_0_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_0_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_0_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_1_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_1_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_1_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_2_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_2_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_2_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_3_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_3_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_3_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_4_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_4_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_4_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_5_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_5_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_5_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_6_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_6_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_6_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_7_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_7_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_7_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_8_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_8_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_8_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_9_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_9_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_9_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_10_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_10_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_10_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_11_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_11_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_11_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_12_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_12_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_12_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_13_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_13_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_13_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_14_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_14_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_14_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_15_ready; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_in_15_valid; // @[BFS.scala 903:46]
  wire [31:0] tier_fifo_1_io_in_15_bits_tdata; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_out_full; // @[BFS.scala 903:46]
  wire [511:0] tier_fifo_1_io_out_din; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_out_wr_en; // @[BFS.scala 903:46]
  wire [511:0] tier_fifo_1_io_out_dout; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_out_rd_en; // @[BFS.scala 903:46]
  wire [8:0] tier_fifo_1_io_out_data_count; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_out_valid; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_flush; // @[BFS.scala 903:46]
  wire  tier_fifo_1_io_is_current_tier; // @[BFS.scala 903:46]
  (*dont_touch = "true" *)reg [31:0] tier_counter_0; // @[BFS.scala 904:29]
  (*dont_touch = "true" *)reg [31:0] tier_counter_1; // @[BFS.scala 904:29]
  reg [4:0] status; // @[BFS.scala 922:23]
  reg [4:0] tier_status_0; // @[BFS.scala 923:28]
  reg [4:0] tier_status_1; // @[BFS.scala 923:28]
  wire  _T_1 = io_start & status == 5'h0; // @[BFS.scala 925:17]
  wire  _T_2 = status == 5'h2; // @[BFS.scala 927:21]
  wire  _T_5 = status == 5'h5; // @[BFS.scala 929:21]
  wire  _T_8 = status == 5'h7; // @[BFS.scala 931:34]
  wire [4:0] _GEN_0 = tier_status_1 != 5'h0 ? 5'h12 : 5'h1; // @[BFS.scala 932:39 BFS.scala 933:14 BFS.scala 935:14]
  wire  _T_11 = status == 5'h1; // @[BFS.scala 937:21]
  wire  _T_14 = status == 5'h6; // @[BFS.scala 939:21]
  wire  _T_17 = status == 5'h8; // @[BFS.scala 941:34]
  wire [4:0] _GEN_1 = tier_status_0 != 5'h0 ? 5'h11 : 5'h2; // @[BFS.scala 942:38 BFS.scala 943:14 BFS.scala 945:14]
  wire  _T_20 = status == 5'h11; // @[BFS.scala 947:21]
  wire  _T_21 = tier_status_0 == 5'h0; // @[BFS.scala 947:60]
  wire  _T_23 = status == 5'h12; // @[BFS.scala 949:21]
  wire  _T_24 = tier_status_1 == 5'h0; // @[BFS.scala 949:60]
  wire [4:0] _GEN_2 = io_end ? 5'h0 : status; // @[BFS.scala 951:21 BFS.scala 952:12 BFS.scala 922:23]
  wire [4:0] _GEN_3 = status == 5'h12 & tier_status_1 == 5'h0 ? 5'h1 : _GEN_2; // @[BFS.scala 949:73 BFS.scala 950:12]
  wire [4:0] _GEN_4 = status == 5'h11 & tier_status_0 == 5'h0 ? 5'h2 : _GEN_3; // @[BFS.scala 947:73 BFS.scala 948:12]
  wire [4:0] _GEN_5 = io_signal & status == 5'h8 ? _GEN_1 : _GEN_4; // @[BFS.scala 941:55]
  wire [4:0] _GEN_6 = status == 5'h6 & io_cacheable_out_valid & io_cacheable_out_ready ? 5'h8 : _GEN_5; // @[BFS.scala 939:92 BFS.scala 940:12]
  wire [4:0] _GEN_7 = status == 5'h1 & tier_counter_1 == 32'h0 ? 5'h6 : _GEN_6; // @[BFS.scala 937:70 BFS.scala 938:12]
  wire [4:0] _GEN_8 = io_signal & status == 5'h7 ? _GEN_0 : _GEN_7; // @[BFS.scala 931:55]
  wire  next_tier_mask_hi = _T_2 | _T_5 | _T_8 | _T_23; // @[BFS.scala 955:115]
  wire  next_tier_mask_lo = _T_11 | _T_14 | _T_17 | _T_20; // @[BFS.scala 956:94]
  wire [1:0] next_tier_mask = {next_tier_mask_hi,next_tier_mask_lo}; // @[Cat.scala 30:58]
  reg [63:0] tier_base_addr_0; // @[BFS.scala 958:31]
  reg [63:0] tier_base_addr_1; // @[BFS.scala 958:31]
  wire  _step_fin_T_2 = _T_8 | _T_17; // @[BFS.scala 959:60]
  wire  step_fin = io_signal & (_T_8 | _T_17); // @[BFS.scala 959:28]
  wire  _axi_aw_valid_T_1 = tier_status_0 == 5'h3; // @[BFS.scala 1045:57]
  wire  _axi_aw_valid_T_2 = tier_status_1 == 5'h3; // @[BFS.scala 1045:90]
  wire  axi_aw_valid = next_tier_mask[0] ? tier_status_0 == 5'h3 : tier_status_1 == 5'h3; // @[BFS.scala 1045:22]
  wire [63:0] _tier_base_addr_0_T_1 = tier_base_addr_0 + 64'h400; // @[BFS.scala 965:16]
  wire  _T_35 = ~next_tier_mask[0]; // @[BFS.scala 966:18]
  wire  _axi_ar_valid_T_1 = tier_status_1 == 5'h4; // @[BFS.scala 1052:57]
  wire  _axi_ar_valid_T_2 = tier_status_0 == 5'h4; // @[BFS.scala 1052:89]
  wire  axi_ar_valid = next_tier_mask[0] ? tier_status_1 == 5'h4 : tier_status_0 == 5'h4; // @[BFS.scala 1052:22]
  wire [63:0] _tier_base_addr_1_T_1 = tier_base_addr_1 + 64'h400; // @[BFS.scala 965:16]
  wire  _T_49 = ~next_tier_mask[1]; // @[BFS.scala 966:18]
  wire  _T_55 = io_cacheable_in_0_ready & io_cacheable_in_0_valid; // @[BFS.scala 973:72]
  wire  _T_56 = io_cacheable_in_1_ready & io_cacheable_in_1_valid; // @[BFS.scala 973:72]
  wire  _T_57 = io_cacheable_in_2_ready & io_cacheable_in_2_valid; // @[BFS.scala 973:72]
  wire  _T_58 = io_cacheable_in_3_ready & io_cacheable_in_3_valid; // @[BFS.scala 973:72]
  wire  _T_59 = io_cacheable_in_4_ready & io_cacheable_in_4_valid; // @[BFS.scala 973:72]
  wire  _T_60 = io_cacheable_in_5_ready & io_cacheable_in_5_valid; // @[BFS.scala 973:72]
  wire  _T_61 = io_cacheable_in_6_ready & io_cacheable_in_6_valid; // @[BFS.scala 973:72]
  wire  _T_62 = io_cacheable_in_7_ready & io_cacheable_in_7_valid; // @[BFS.scala 973:72]
  wire  _T_63 = io_cacheable_in_8_ready & io_cacheable_in_8_valid; // @[BFS.scala 973:72]
  wire  _T_64 = io_cacheable_in_9_ready & io_cacheable_in_9_valid; // @[BFS.scala 973:72]
  wire  _T_65 = io_cacheable_in_10_ready & io_cacheable_in_10_valid; // @[BFS.scala 973:72]
  wire  _T_66 = io_cacheable_in_11_ready & io_cacheable_in_11_valid; // @[BFS.scala 973:72]
  wire  _T_67 = io_cacheable_in_12_ready & io_cacheable_in_12_valid; // @[BFS.scala 973:72]
  wire  _T_68 = io_cacheable_in_13_ready & io_cacheable_in_13_valid; // @[BFS.scala 973:72]
  wire  _T_69 = io_cacheable_in_14_ready & io_cacheable_in_14_valid; // @[BFS.scala 973:72]
  wire  _T_70 = io_cacheable_in_15_ready & io_cacheable_in_15_valid; // @[BFS.scala 973:72]
  wire  _T_85 = io_cacheable_in_0_ready & io_cacheable_in_0_valid | io_cacheable_in_1_ready & io_cacheable_in_1_valid |
    io_cacheable_in_2_ready & io_cacheable_in_2_valid | io_cacheable_in_3_ready & io_cacheable_in_3_valid |
    io_cacheable_in_4_ready & io_cacheable_in_4_valid | io_cacheable_in_5_ready & io_cacheable_in_5_valid |
    io_cacheable_in_6_ready & io_cacheable_in_6_valid | io_cacheable_in_7_ready & io_cacheable_in_7_valid |
    io_cacheable_in_8_ready & io_cacheable_in_8_valid | io_cacheable_in_9_ready & io_cacheable_in_9_valid |
    io_cacheable_in_10_ready & io_cacheable_in_10_valid | io_cacheable_in_11_ready & io_cacheable_in_11_valid |
    io_cacheable_in_12_ready & io_cacheable_in_12_valid | io_cacheable_in_13_ready & io_cacheable_in_13_valid |
    io_cacheable_in_14_ready & io_cacheable_in_14_valid | _T_70; // @[BFS.scala 973:93]
  wire [5:0] _tier_counter_0_WIRE = {{5'd0}, _T_55}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_WIRE_1 = {{5'd0}, _T_56}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_17 = _tier_counter_0_WIRE + _tier_counter_0_WIRE_1; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_2 = {{5'd0}, _T_57}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_19 = _tier_counter_0_T_17 + _tier_counter_0_WIRE_2; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_3 = {{5'd0}, _T_58}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_21 = _tier_counter_0_T_19 + _tier_counter_0_WIRE_3; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_4 = {{5'd0}, _T_59}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_23 = _tier_counter_0_T_21 + _tier_counter_0_WIRE_4; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_5 = {{5'd0}, _T_60}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_25 = _tier_counter_0_T_23 + _tier_counter_0_WIRE_5; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_6 = {{5'd0}, _T_61}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_27 = _tier_counter_0_T_25 + _tier_counter_0_WIRE_6; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_7 = {{5'd0}, _T_62}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_29 = _tier_counter_0_T_27 + _tier_counter_0_WIRE_7; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_8 = {{5'd0}, _T_63}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_31 = _tier_counter_0_T_29 + _tier_counter_0_WIRE_8; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_9 = {{5'd0}, _T_64}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_33 = _tier_counter_0_T_31 + _tier_counter_0_WIRE_9; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_10 = {{5'd0}, _T_65}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_35 = _tier_counter_0_T_33 + _tier_counter_0_WIRE_10; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_11 = {{5'd0}, _T_66}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_37 = _tier_counter_0_T_35 + _tier_counter_0_WIRE_11; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_12 = {{5'd0}, _T_67}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_39 = _tier_counter_0_T_37 + _tier_counter_0_WIRE_12; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_13 = {{5'd0}, _T_68}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_41 = _tier_counter_0_T_39 + _tier_counter_0_WIRE_13; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_14 = {{5'd0}, _T_69}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_43 = _tier_counter_0_T_41 + _tier_counter_0_WIRE_14; // @[BFS.scala 974:100]
  wire [5:0] _tier_counter_0_WIRE_15 = {{5'd0}, _T_70}; // @[BFS.scala 974:78 BFS.scala 974:78]
  wire [5:0] _tier_counter_0_T_45 = _tier_counter_0_T_43 + _tier_counter_0_WIRE_15; // @[BFS.scala 974:100]
  wire [31:0] _GEN_36 = {{26'd0}, _tier_counter_0_T_45}; // @[BFS.scala 974:16]
  wire [31:0] _tier_counter_0_T_47 = tier_counter_0 + _GEN_36; // @[BFS.scala 974:16]
  wire [31:0] _tier_counter_0_T_50 = tier_counter_0 - 32'h10; // @[BFS.scala 976:59]
  wire [31:0] _GEN_37 = {{23'd0}, tier_fifo_0_io_out_data_count}; // @[BFS.scala 976:69]
  wire [31:0] _tier_counter_0_T_52 = tier_counter_0 - _GEN_37; // @[BFS.scala 976:69]
  wire [31:0] _tier_counter_1_T_47 = tier_counter_1 + _GEN_36; // @[BFS.scala 974:16]
  wire [31:0] _tier_counter_1_T_50 = tier_counter_1 - 32'h10; // @[BFS.scala 976:59]
  wire [31:0] _GEN_39 = {{23'd0}, tier_fifo_1_io_out_data_count}; // @[BFS.scala 976:69]
  wire [31:0] _tier_counter_1_T_52 = tier_counter_1 - _GEN_39; // @[BFS.scala 976:69]
  wire  _T_134 = tier_fifo_0_io_out_data_count == 9'h0; // @[BFS.scala 818:23]
  wire  _T_149 = tier_status_0 == 5'h9; // @[BFS.scala 1007:20]
  reg [7:0] wcount; // @[BFS.scala 1033:23]
  wire  axi_w_bits_wlast = wcount == 8'h1; // @[BFS.scala 1055:30]
  wire [4:0] _GEN_22 = tier_status_0 == 5'h9 & axi_w_bits_wlast & io_ddr_out_0_w_ready ? 5'h0 : tier_status_0; // @[BFS.scala 1007:94 BFS.scala 1008:11 BFS.scala 923:28]
  wire [4:0] _GEN_23 = tier_status_0 == 5'h10 & io_ddr_out_0_r_bits_rlast & io_ddr_out_0_r_valid ? 5'h0 : _GEN_22; // @[BFS.scala 1005:99 BFS.scala 1006:11]
  wire [4:0] _GEN_24 = _axi_ar_valid_T_2 & io_ddr_out_0_ar_ready ? 5'h10 : _GEN_23; // @[BFS.scala 1003:52 BFS.scala 1004:11]
  wire  _T_160 = tier_fifo_1_io_out_data_count == 9'h0; // @[BFS.scala 818:23]
  wire  _T_175 = tier_status_1 == 5'h9; // @[BFS.scala 1007:20]
  wire [4:0] _GEN_28 = tier_status_1 == 5'h9 & axi_w_bits_wlast & io_ddr_out_0_w_ready ? 5'h0 : tier_status_1; // @[BFS.scala 1007:94 BFS.scala 1008:11 BFS.scala 923:28]
  wire [4:0] _GEN_29 = tier_status_1 == 5'h10 & io_ddr_out_0_r_bits_rlast & io_ddr_out_0_r_valid ? 5'h0 : _GEN_28; // @[BFS.scala 1005:99 BFS.scala 1006:11]
  wire [4:0] _GEN_30 = _axi_ar_valid_T_1 & io_ddr_out_0_ar_ready ? 5'h10 : _GEN_29; // @[BFS.scala 1003:52 BFS.scala 1004:11]
  wire  _io_cacheable_out_valid_T_2 = tier_fifo_1_io_out_valid | _T_14; // @[BFS.scala 1020:57]
  wire  _io_cacheable_out_valid_T_5 = tier_fifo_0_io_out_valid | _T_5; // @[BFS.scala 1021:57]
  wire [511:0] _io_cacheable_out_bits_tdata_T_4 = next_tier_mask[1] ? tier_fifo_0_io_out_dout : 512'h0; // @[Mux.scala 98:16]
  wire [511:0] _io_cacheable_out_bits_tdata_T_5 = next_tier_mask[0] ? tier_fifo_1_io_out_dout :
    _io_cacheable_out_bits_tdata_T_4; // @[Mux.scala 98:16]
  wire [511:0] _io_cacheable_out_bits_tdata_T_6 = _T_14 ? 512'h80000000 : _io_cacheable_out_bits_tdata_T_5; // @[Mux.scala 98:16]
  wire  _io_cacheable_out_bits_tkeep_T_6 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h0 :
    tier_fifo_0_io_out_data_count > 9'h0; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_10 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h1 :
    tier_fifo_0_io_out_data_count > 9'h1; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_14 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h2 :
    tier_fifo_0_io_out_data_count > 9'h2; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_18 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h3 :
    tier_fifo_0_io_out_data_count > 9'h3; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_22 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h4 :
    tier_fifo_0_io_out_data_count > 9'h4; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_26 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h5 :
    tier_fifo_0_io_out_data_count > 9'h5; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_30 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h6 :
    tier_fifo_0_io_out_data_count > 9'h6; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_34 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h7 :
    tier_fifo_0_io_out_data_count > 9'h7; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_38 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h8 :
    tier_fifo_0_io_out_data_count > 9'h8; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_42 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'h9 :
    tier_fifo_0_io_out_data_count > 9'h9; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_46 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'ha :
    tier_fifo_0_io_out_data_count > 9'ha; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_50 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'hb :
    tier_fifo_0_io_out_data_count > 9'hb; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_54 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'hc :
    tier_fifo_0_io_out_data_count > 9'hc; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_58 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'hd :
    tier_fifo_0_io_out_data_count > 9'hd; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_62 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'he :
    tier_fifo_0_io_out_data_count > 9'he; // @[BFS.scala 1029:15]
  wire  _io_cacheable_out_bits_tkeep_T_66 = next_tier_mask[0] ? tier_fifo_1_io_out_data_count > 9'hf :
    tier_fifo_0_io_out_data_count > 9'hf; // @[BFS.scala 1029:15]
  wire [7:0] io_cacheable_out_bits_tkeep_lo = {_io_cacheable_out_bits_tkeep_T_34,_io_cacheable_out_bits_tkeep_T_30,
    _io_cacheable_out_bits_tkeep_T_26,_io_cacheable_out_bits_tkeep_T_22,_io_cacheable_out_bits_tkeep_T_18,
    _io_cacheable_out_bits_tkeep_T_14,_io_cacheable_out_bits_tkeep_T_10,_io_cacheable_out_bits_tkeep_T_6}; // @[BFS.scala 1030:14]
  wire [15:0] _io_cacheable_out_bits_tkeep_T_67 = {_io_cacheable_out_bits_tkeep_T_66,_io_cacheable_out_bits_tkeep_T_62,
    _io_cacheable_out_bits_tkeep_T_58,_io_cacheable_out_bits_tkeep_T_54,_io_cacheable_out_bits_tkeep_T_50,
    _io_cacheable_out_bits_tkeep_T_46,_io_cacheable_out_bits_tkeep_T_42,_io_cacheable_out_bits_tkeep_T_38,
    io_cacheable_out_bits_tkeep_lo}; // @[BFS.scala 1030:14]
  wire  axi_w_valid = next_tier_mask[0] ? _T_149 : _T_175; // @[BFS.scala 1054:21]
  wire [7:0] _wcount_T_1 = wcount - 8'h1; // @[BFS.scala 1037:22]
  multi_channel_fifo tier_fifo_0 ( // @[BFS.scala 903:46]
    .clock(tier_fifo_0_clock),
    .reset(tier_fifo_0_reset),
    .io_in_0_ready(tier_fifo_0_io_in_0_ready),
    .io_in_0_valid(tier_fifo_0_io_in_0_valid),
    .io_in_0_bits_tdata(tier_fifo_0_io_in_0_bits_tdata),
    .io_in_1_ready(tier_fifo_0_io_in_1_ready),
    .io_in_1_valid(tier_fifo_0_io_in_1_valid),
    .io_in_1_bits_tdata(tier_fifo_0_io_in_1_bits_tdata),
    .io_in_2_ready(tier_fifo_0_io_in_2_ready),
    .io_in_2_valid(tier_fifo_0_io_in_2_valid),
    .io_in_2_bits_tdata(tier_fifo_0_io_in_2_bits_tdata),
    .io_in_3_ready(tier_fifo_0_io_in_3_ready),
    .io_in_3_valid(tier_fifo_0_io_in_3_valid),
    .io_in_3_bits_tdata(tier_fifo_0_io_in_3_bits_tdata),
    .io_in_4_ready(tier_fifo_0_io_in_4_ready),
    .io_in_4_valid(tier_fifo_0_io_in_4_valid),
    .io_in_4_bits_tdata(tier_fifo_0_io_in_4_bits_tdata),
    .io_in_5_ready(tier_fifo_0_io_in_5_ready),
    .io_in_5_valid(tier_fifo_0_io_in_5_valid),
    .io_in_5_bits_tdata(tier_fifo_0_io_in_5_bits_tdata),
    .io_in_6_ready(tier_fifo_0_io_in_6_ready),
    .io_in_6_valid(tier_fifo_0_io_in_6_valid),
    .io_in_6_bits_tdata(tier_fifo_0_io_in_6_bits_tdata),
    .io_in_7_ready(tier_fifo_0_io_in_7_ready),
    .io_in_7_valid(tier_fifo_0_io_in_7_valid),
    .io_in_7_bits_tdata(tier_fifo_0_io_in_7_bits_tdata),
    .io_in_8_ready(tier_fifo_0_io_in_8_ready),
    .io_in_8_valid(tier_fifo_0_io_in_8_valid),
    .io_in_8_bits_tdata(tier_fifo_0_io_in_8_bits_tdata),
    .io_in_9_ready(tier_fifo_0_io_in_9_ready),
    .io_in_9_valid(tier_fifo_0_io_in_9_valid),
    .io_in_9_bits_tdata(tier_fifo_0_io_in_9_bits_tdata),
    .io_in_10_ready(tier_fifo_0_io_in_10_ready),
    .io_in_10_valid(tier_fifo_0_io_in_10_valid),
    .io_in_10_bits_tdata(tier_fifo_0_io_in_10_bits_tdata),
    .io_in_11_ready(tier_fifo_0_io_in_11_ready),
    .io_in_11_valid(tier_fifo_0_io_in_11_valid),
    .io_in_11_bits_tdata(tier_fifo_0_io_in_11_bits_tdata),
    .io_in_12_ready(tier_fifo_0_io_in_12_ready),
    .io_in_12_valid(tier_fifo_0_io_in_12_valid),
    .io_in_12_bits_tdata(tier_fifo_0_io_in_12_bits_tdata),
    .io_in_13_ready(tier_fifo_0_io_in_13_ready),
    .io_in_13_valid(tier_fifo_0_io_in_13_valid),
    .io_in_13_bits_tdata(tier_fifo_0_io_in_13_bits_tdata),
    .io_in_14_ready(tier_fifo_0_io_in_14_ready),
    .io_in_14_valid(tier_fifo_0_io_in_14_valid),
    .io_in_14_bits_tdata(tier_fifo_0_io_in_14_bits_tdata),
    .io_in_15_ready(tier_fifo_0_io_in_15_ready),
    .io_in_15_valid(tier_fifo_0_io_in_15_valid),
    .io_in_15_bits_tdata(tier_fifo_0_io_in_15_bits_tdata),
    .io_out_full(tier_fifo_0_io_out_full),
    .io_out_din(tier_fifo_0_io_out_din),
    .io_out_wr_en(tier_fifo_0_io_out_wr_en),
    .io_out_dout(tier_fifo_0_io_out_dout),
    .io_out_rd_en(tier_fifo_0_io_out_rd_en),
    .io_out_data_count(tier_fifo_0_io_out_data_count),
    .io_out_valid(tier_fifo_0_io_out_valid),
    .io_flush(tier_fifo_0_io_flush),
    .io_is_current_tier(tier_fifo_0_io_is_current_tier)
  );
  multi_channel_fifo tier_fifo_1 ( // @[BFS.scala 903:46]
    .clock(tier_fifo_1_clock),
    .reset(tier_fifo_1_reset),
    .io_in_0_ready(tier_fifo_1_io_in_0_ready),
    .io_in_0_valid(tier_fifo_1_io_in_0_valid),
    .io_in_0_bits_tdata(tier_fifo_1_io_in_0_bits_tdata),
    .io_in_1_ready(tier_fifo_1_io_in_1_ready),
    .io_in_1_valid(tier_fifo_1_io_in_1_valid),
    .io_in_1_bits_tdata(tier_fifo_1_io_in_1_bits_tdata),
    .io_in_2_ready(tier_fifo_1_io_in_2_ready),
    .io_in_2_valid(tier_fifo_1_io_in_2_valid),
    .io_in_2_bits_tdata(tier_fifo_1_io_in_2_bits_tdata),
    .io_in_3_ready(tier_fifo_1_io_in_3_ready),
    .io_in_3_valid(tier_fifo_1_io_in_3_valid),
    .io_in_3_bits_tdata(tier_fifo_1_io_in_3_bits_tdata),
    .io_in_4_ready(tier_fifo_1_io_in_4_ready),
    .io_in_4_valid(tier_fifo_1_io_in_4_valid),
    .io_in_4_bits_tdata(tier_fifo_1_io_in_4_bits_tdata),
    .io_in_5_ready(tier_fifo_1_io_in_5_ready),
    .io_in_5_valid(tier_fifo_1_io_in_5_valid),
    .io_in_5_bits_tdata(tier_fifo_1_io_in_5_bits_tdata),
    .io_in_6_ready(tier_fifo_1_io_in_6_ready),
    .io_in_6_valid(tier_fifo_1_io_in_6_valid),
    .io_in_6_bits_tdata(tier_fifo_1_io_in_6_bits_tdata),
    .io_in_7_ready(tier_fifo_1_io_in_7_ready),
    .io_in_7_valid(tier_fifo_1_io_in_7_valid),
    .io_in_7_bits_tdata(tier_fifo_1_io_in_7_bits_tdata),
    .io_in_8_ready(tier_fifo_1_io_in_8_ready),
    .io_in_8_valid(tier_fifo_1_io_in_8_valid),
    .io_in_8_bits_tdata(tier_fifo_1_io_in_8_bits_tdata),
    .io_in_9_ready(tier_fifo_1_io_in_9_ready),
    .io_in_9_valid(tier_fifo_1_io_in_9_valid),
    .io_in_9_bits_tdata(tier_fifo_1_io_in_9_bits_tdata),
    .io_in_10_ready(tier_fifo_1_io_in_10_ready),
    .io_in_10_valid(tier_fifo_1_io_in_10_valid),
    .io_in_10_bits_tdata(tier_fifo_1_io_in_10_bits_tdata),
    .io_in_11_ready(tier_fifo_1_io_in_11_ready),
    .io_in_11_valid(tier_fifo_1_io_in_11_valid),
    .io_in_11_bits_tdata(tier_fifo_1_io_in_11_bits_tdata),
    .io_in_12_ready(tier_fifo_1_io_in_12_ready),
    .io_in_12_valid(tier_fifo_1_io_in_12_valid),
    .io_in_12_bits_tdata(tier_fifo_1_io_in_12_bits_tdata),
    .io_in_13_ready(tier_fifo_1_io_in_13_ready),
    .io_in_13_valid(tier_fifo_1_io_in_13_valid),
    .io_in_13_bits_tdata(tier_fifo_1_io_in_13_bits_tdata),
    .io_in_14_ready(tier_fifo_1_io_in_14_ready),
    .io_in_14_valid(tier_fifo_1_io_in_14_valid),
    .io_in_14_bits_tdata(tier_fifo_1_io_in_14_bits_tdata),
    .io_in_15_ready(tier_fifo_1_io_in_15_ready),
    .io_in_15_valid(tier_fifo_1_io_in_15_valid),
    .io_in_15_bits_tdata(tier_fifo_1_io_in_15_bits_tdata),
    .io_out_full(tier_fifo_1_io_out_full),
    .io_out_din(tier_fifo_1_io_out_din),
    .io_out_wr_en(tier_fifo_1_io_out_wr_en),
    .io_out_dout(tier_fifo_1_io_out_dout),
    .io_out_rd_en(tier_fifo_1_io_out_rd_en),
    .io_out_data_count(tier_fifo_1_io_out_data_count),
    .io_out_valid(tier_fifo_1_io_out_valid),
    .io_flush(tier_fifo_1_io_flush),
    .io_is_current_tier(tier_fifo_1_io_is_current_tier)
  );
  assign io_cacheable_out_valid = next_tier_mask[0] ? _io_cacheable_out_valid_T_2 : next_tier_mask[1] &
    _io_cacheable_out_valid_T_5; // @[Mux.scala 98:16]
  assign io_cacheable_out_bits_tdata = _T_5 ? 512'h80000000 : _io_cacheable_out_bits_tdata_T_6; // @[Mux.scala 98:16]
  assign io_cacheable_out_bits_tkeep = _T_5 | _T_14 ? 16'h1 : _io_cacheable_out_bits_tkeep_T_67; // @[BFS.scala 1027:37]
  assign io_cacheable_in_0_ready = next_tier_mask[0] ? tier_fifo_0_io_in_0_ready : tier_fifo_1_io_in_0_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_1_ready = next_tier_mask[0] ? tier_fifo_0_io_in_1_ready : tier_fifo_1_io_in_1_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_2_ready = next_tier_mask[0] ? tier_fifo_0_io_in_2_ready : tier_fifo_1_io_in_2_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_3_ready = next_tier_mask[0] ? tier_fifo_0_io_in_3_ready : tier_fifo_1_io_in_3_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_4_ready = next_tier_mask[0] ? tier_fifo_0_io_in_4_ready : tier_fifo_1_io_in_4_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_5_ready = next_tier_mask[0] ? tier_fifo_0_io_in_5_ready : tier_fifo_1_io_in_5_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_6_ready = next_tier_mask[0] ? tier_fifo_0_io_in_6_ready : tier_fifo_1_io_in_6_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_7_ready = next_tier_mask[0] ? tier_fifo_0_io_in_7_ready : tier_fifo_1_io_in_7_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_8_ready = next_tier_mask[0] ? tier_fifo_0_io_in_8_ready : tier_fifo_1_io_in_8_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_9_ready = next_tier_mask[0] ? tier_fifo_0_io_in_9_ready : tier_fifo_1_io_in_9_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_10_ready = next_tier_mask[0] ? tier_fifo_0_io_in_10_ready : tier_fifo_1_io_in_10_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_11_ready = next_tier_mask[0] ? tier_fifo_0_io_in_11_ready : tier_fifo_1_io_in_11_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_12_ready = next_tier_mask[0] ? tier_fifo_0_io_in_12_ready : tier_fifo_1_io_in_12_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_13_ready = next_tier_mask[0] ? tier_fifo_0_io_in_13_ready : tier_fifo_1_io_in_13_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_14_ready = next_tier_mask[0] ? tier_fifo_0_io_in_14_ready : tier_fifo_1_io_in_14_ready; // @[BFS.scala 1015:22]
  assign io_cacheable_in_15_ready = next_tier_mask[0] ? tier_fifo_0_io_in_15_ready : tier_fifo_1_io_in_15_ready; // @[BFS.scala 1015:22]
  assign io_non_cacheable_in_aw_ready = io_ddr_out_1_aw_ready; // @[BFS.scala 1061:17]
  assign io_non_cacheable_in_w_ready = io_ddr_out_1_w_ready; // @[BFS.scala 1061:17]
  assign io_ddr_out_0_aw_valid = next_tier_mask[0] ? tier_status_0 == 5'h3 : tier_status_1 == 5'h3; // @[BFS.scala 1045:22]
  assign io_ddr_out_0_aw_bits_awaddr = next_tier_mask[0] ? tier_base_addr_0 : tier_base_addr_1; // @[BFS.scala 1039:28]
  assign io_ddr_out_0_ar_valid = next_tier_mask[0] ? tier_status_1 == 5'h4 : tier_status_0 == 5'h4; // @[BFS.scala 1052:22]
  assign io_ddr_out_0_ar_bits_araddr = next_tier_mask[0] ? tier_base_addr_1 : tier_base_addr_0; // @[BFS.scala 1046:28]
  assign io_ddr_out_0_w_valid = next_tier_mask[0] ? _T_149 : _T_175; // @[BFS.scala 1054:21]
  assign io_ddr_out_0_w_bits_wdata = next_tier_mask[0] ? tier_fifo_0_io_out_dout : tier_fifo_1_io_out_dout; // @[BFS.scala 1053:26]
  assign io_ddr_out_0_w_bits_wlast = wcount == 8'h1; // @[BFS.scala 1055:30]
  assign io_ddr_out_1_aw_valid = io_non_cacheable_in_aw_valid; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_aw_bits_awaddr = io_non_cacheable_in_aw_bits_awaddr; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_aw_bits_awid = io_non_cacheable_in_aw_bits_awid; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_w_valid = io_non_cacheable_in_w_valid; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_w_bits_wdata = io_non_cacheable_in_w_bits_wdata; // @[BFS.scala 1061:17]
  assign io_ddr_out_1_w_bits_wstrb = io_non_cacheable_in_w_bits_wstrb; // @[BFS.scala 1061:17]
  assign io_unvisited_size = next_tier_mask[0] ? tier_counter_0 : tier_counter_1; // @[BFS.scala 1018:27]
  assign io_signal_ack = _T_17 | _T_8; // @[BFS.scala 1063:48]
  assign tier_fifo_0_clock = clock;
  assign tier_fifo_0_reset = reset;
  assign tier_fifo_0_io_in_0_valid = next_tier_mask[0] & io_cacheable_in_0_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_0_bits_tdata = next_tier_mask[0] ? io_cacheable_in_0_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_1_valid = next_tier_mask[0] & io_cacheable_in_1_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_1_bits_tdata = next_tier_mask[0] ? io_cacheable_in_1_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_2_valid = next_tier_mask[0] & io_cacheable_in_2_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_2_bits_tdata = next_tier_mask[0] ? io_cacheable_in_2_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_3_valid = next_tier_mask[0] & io_cacheable_in_3_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_3_bits_tdata = next_tier_mask[0] ? io_cacheable_in_3_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_4_valid = next_tier_mask[0] & io_cacheable_in_4_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_4_bits_tdata = next_tier_mask[0] ? io_cacheable_in_4_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_5_valid = next_tier_mask[0] & io_cacheable_in_5_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_5_bits_tdata = next_tier_mask[0] ? io_cacheable_in_5_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_6_valid = next_tier_mask[0] & io_cacheable_in_6_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_6_bits_tdata = next_tier_mask[0] ? io_cacheable_in_6_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_7_valid = next_tier_mask[0] & io_cacheable_in_7_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_7_bits_tdata = next_tier_mask[0] ? io_cacheable_in_7_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_8_valid = next_tier_mask[0] & io_cacheable_in_8_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_8_bits_tdata = next_tier_mask[0] ? io_cacheable_in_8_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_9_valid = next_tier_mask[0] & io_cacheable_in_9_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_9_bits_tdata = next_tier_mask[0] ? io_cacheable_in_9_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_10_valid = next_tier_mask[0] & io_cacheable_in_10_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_10_bits_tdata = next_tier_mask[0] ? io_cacheable_in_10_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_11_valid = next_tier_mask[0] & io_cacheable_in_11_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_11_bits_tdata = next_tier_mask[0] ? io_cacheable_in_11_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_12_valid = next_tier_mask[0] & io_cacheable_in_12_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_12_bits_tdata = next_tier_mask[0] ? io_cacheable_in_12_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_13_valid = next_tier_mask[0] & io_cacheable_in_13_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_13_bits_tdata = next_tier_mask[0] ? io_cacheable_in_13_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_14_valid = next_tier_mask[0] & io_cacheable_in_14_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_14_bits_tdata = next_tier_mask[0] ? io_cacheable_in_14_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_in_15_valid = next_tier_mask[0] & io_cacheable_in_15_valid; // @[BFS.scala 988:26]
  assign tier_fifo_0_io_in_15_bits_tdata = next_tier_mask[0] ? io_cacheable_in_15_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_0_io_out_din = next_tier_mask[0] ? 512'h0 : io_ddr_out_0_r_bits_rdata; // @[BFS.scala 984:26]
  assign tier_fifo_0_io_out_wr_en = next_tier_mask[0] ? 1'h0 : io_ddr_out_0_r_valid; // @[BFS.scala 983:28]
  assign tier_fifo_0_io_out_rd_en = next_tier_mask[0] ? io_ddr_out_0_w_ready : io_cacheable_out_ready; // @[BFS.scala 982:28]
  assign tier_fifo_0_io_flush = io_signal & _step_fin_T_2; // @[BFS.scala 985:31]
  assign tier_fifo_0_io_is_current_tier = ~next_tier_mask[0]; // @[BFS.scala 992:31]
  assign tier_fifo_1_clock = clock;
  assign tier_fifo_1_reset = reset;
  assign tier_fifo_1_io_in_0_valid = next_tier_mask[1] & io_cacheable_in_0_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_0_bits_tdata = next_tier_mask[1] ? io_cacheable_in_0_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_1_valid = next_tier_mask[1] & io_cacheable_in_1_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_1_bits_tdata = next_tier_mask[1] ? io_cacheable_in_1_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_2_valid = next_tier_mask[1] & io_cacheable_in_2_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_2_bits_tdata = next_tier_mask[1] ? io_cacheable_in_2_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_3_valid = next_tier_mask[1] & io_cacheable_in_3_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_3_bits_tdata = next_tier_mask[1] ? io_cacheable_in_3_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_4_valid = next_tier_mask[1] & io_cacheable_in_4_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_4_bits_tdata = next_tier_mask[1] ? io_cacheable_in_4_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_5_valid = next_tier_mask[1] & io_cacheable_in_5_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_5_bits_tdata = next_tier_mask[1] ? io_cacheable_in_5_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_6_valid = next_tier_mask[1] & io_cacheable_in_6_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_6_bits_tdata = next_tier_mask[1] ? io_cacheable_in_6_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_7_valid = next_tier_mask[1] & io_cacheable_in_7_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_7_bits_tdata = next_tier_mask[1] ? io_cacheable_in_7_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_8_valid = next_tier_mask[1] & io_cacheable_in_8_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_8_bits_tdata = next_tier_mask[1] ? io_cacheable_in_8_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_9_valid = next_tier_mask[1] & io_cacheable_in_9_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_9_bits_tdata = next_tier_mask[1] ? io_cacheable_in_9_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_10_valid = next_tier_mask[1] & io_cacheable_in_10_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_10_bits_tdata = next_tier_mask[1] ? io_cacheable_in_10_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_11_valid = next_tier_mask[1] & io_cacheable_in_11_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_11_bits_tdata = next_tier_mask[1] ? io_cacheable_in_11_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_12_valid = next_tier_mask[1] & io_cacheable_in_12_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_12_bits_tdata = next_tier_mask[1] ? io_cacheable_in_12_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_13_valid = next_tier_mask[1] & io_cacheable_in_13_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_13_bits_tdata = next_tier_mask[1] ? io_cacheable_in_13_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_14_valid = next_tier_mask[1] & io_cacheable_in_14_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_14_bits_tdata = next_tier_mask[1] ? io_cacheable_in_14_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_in_15_valid = next_tier_mask[1] & io_cacheable_in_15_valid; // @[BFS.scala 988:26]
  assign tier_fifo_1_io_in_15_bits_tdata = next_tier_mask[1] ? io_cacheable_in_15_bits_tdata : 32'h0; // @[BFS.scala 989:25]
  assign tier_fifo_1_io_out_din = next_tier_mask[1] ? 512'h0 : io_ddr_out_0_r_bits_rdata; // @[BFS.scala 984:26]
  assign tier_fifo_1_io_out_wr_en = next_tier_mask[1] ? 1'h0 : io_ddr_out_0_r_valid; // @[BFS.scala 983:28]
  assign tier_fifo_1_io_out_rd_en = next_tier_mask[1] ? io_ddr_out_0_w_ready : io_cacheable_out_ready; // @[BFS.scala 982:28]
  assign tier_fifo_1_io_flush = io_signal & _step_fin_T_2; // @[BFS.scala 985:31]
  assign tier_fifo_1_io_is_current_tier = ~next_tier_mask[1]; // @[BFS.scala 992:31]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 904:29]
      tier_counter_0 <= 32'h0; // @[BFS.scala 904:29]
    end else if (next_tier_mask[0] & _T_85) begin // @[BFS.scala 973:97]
      tier_counter_0 <= _tier_counter_0_T_47; // @[BFS.scala 974:11]
    end else if (_T_35 & io_cacheable_out_ready & io_cacheable_out_valid) begin // @[BFS.scala 975:89]
      if (tier_fifo_0_io_out_data_count > 9'h10) begin // @[BFS.scala 976:17]
        tier_counter_0 <= _tier_counter_0_T_50;
      end else begin
        tier_counter_0 <= _tier_counter_0_T_52;
      end
    end
    if (reset) begin // @[BFS.scala 904:29]
      tier_counter_1 <= 32'h0; // @[BFS.scala 904:29]
    end else if (next_tier_mask[1] & _T_85) begin // @[BFS.scala 973:97]
      tier_counter_1 <= _tier_counter_1_T_47; // @[BFS.scala 974:11]
    end else if (_T_49 & io_cacheable_out_ready & io_cacheable_out_valid) begin // @[BFS.scala 975:89]
      if (tier_fifo_1_io_out_data_count > 9'h10) begin // @[BFS.scala 976:17]
        tier_counter_1 <= _tier_counter_1_T_50;
      end else begin
        tier_counter_1 <= _tier_counter_1_T_52;
      end
    end
    if (reset) begin // @[BFS.scala 922:23]
      status <= 5'h0; // @[BFS.scala 922:23]
    end else if (io_start & status == 5'h0) begin // @[BFS.scala 925:40]
      status <= 5'h2; // @[BFS.scala 926:12]
    end else if (status == 5'h2 & tier_counter_0 == 32'h0) begin // @[BFS.scala 927:70]
      status <= 5'h5; // @[BFS.scala 928:12]
    end else if (status == 5'h5 & io_cacheable_out_valid & io_cacheable_out_ready) begin // @[BFS.scala 929:92]
      status <= 5'h7; // @[BFS.scala 930:12]
    end else begin
      status <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 923:28]
      tier_status_0 <= 5'h0; // @[BFS.scala 923:28]
    end else if (next_tier_mask[0] & tier_fifo_0_io_out_full & _T_21) begin // @[BFS.scala 997:76]
      tier_status_0 <= 5'h3; // @[BFS.scala 998:11]
    end else if (_T_35 & _T_134 & tier_counter_0 != 32'h0 & _T_21) begin // @[BFS.scala 999:109]
      tier_status_0 <= 5'h4; // @[BFS.scala 1000:11]
    end else if (_axi_aw_valid_T_1 & io_ddr_out_0_aw_ready) begin // @[BFS.scala 1001:53]
      tier_status_0 <= 5'h9; // @[BFS.scala 1002:11]
    end else begin
      tier_status_0 <= _GEN_24;
    end
    if (reset) begin // @[BFS.scala 923:28]
      tier_status_1 <= 5'h0; // @[BFS.scala 923:28]
    end else if (next_tier_mask[1] & tier_fifo_1_io_out_full & _T_24) begin // @[BFS.scala 997:76]
      tier_status_1 <= 5'h3; // @[BFS.scala 998:11]
    end else if (_T_49 & _T_160 & tier_counter_1 != 32'h0 & _T_24) begin // @[BFS.scala 999:109]
      tier_status_1 <= 5'h4; // @[BFS.scala 1000:11]
    end else if (_axi_aw_valid_T_2 & io_ddr_out_0_aw_ready) begin // @[BFS.scala 1001:53]
      tier_status_1 <= 5'h9; // @[BFS.scala 1002:11]
    end else begin
      tier_status_1 <= _GEN_30;
    end
    if (reset) begin // @[BFS.scala 958:31]
      tier_base_addr_0 <= 64'h0; // @[BFS.scala 958:31]
    end else if (_T_1 | step_fin) begin // @[BFS.scala 962:57]
      tier_base_addr_0 <= io_tiers_base_addr_0; // @[BFS.scala 963:11]
    end else if (next_tier_mask[0] & io_ddr_out_0_aw_ready & axi_aw_valid) begin // @[BFS.scala 964:86]
      tier_base_addr_0 <= _tier_base_addr_0_T_1; // @[BFS.scala 965:11]
    end else if (~next_tier_mask[0] & io_ddr_out_0_ar_ready & axi_ar_valid) begin // @[BFS.scala 966:87]
      tier_base_addr_0 <= _tier_base_addr_0_T_1; // @[BFS.scala 967:11]
    end
    if (reset) begin // @[BFS.scala 958:31]
      tier_base_addr_1 <= 64'h0; // @[BFS.scala 958:31]
    end else if (_T_1 | step_fin) begin // @[BFS.scala 962:57]
      tier_base_addr_1 <= io_tiers_base_addr_1; // @[BFS.scala 963:11]
    end else if (next_tier_mask[1] & io_ddr_out_0_aw_ready & axi_aw_valid) begin // @[BFS.scala 964:86]
      tier_base_addr_1 <= _tier_base_addr_1_T_1; // @[BFS.scala 965:11]
    end else if (~next_tier_mask[1] & io_ddr_out_0_ar_ready & axi_ar_valid) begin // @[BFS.scala 966:87]
      tier_base_addr_1 <= _tier_base_addr_1_T_1; // @[BFS.scala 967:11]
    end
    if (reset) begin // @[BFS.scala 1033:23]
      wcount <= 8'h0; // @[BFS.scala 1033:23]
    end else if (axi_aw_valid & io_ddr_out_0_aw_ready) begin // @[BFS.scala 1034:55]
      wcount <= 8'h10; // @[BFS.scala 1035:12]
    end else if (axi_w_valid & io_ddr_out_0_w_ready) begin // @[BFS.scala 1036:59]
      wcount <= _wcount_T_1; // @[BFS.scala 1037:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tier_counter_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  tier_counter_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  status = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  tier_status_0 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  tier_status_1 = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  tier_base_addr_0 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  tier_base_addr_1 = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  wcount = _RAND_7[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_arbitrator(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [1023:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1023:0] data; // @[BFS.scala 241:21]
  reg [31:0] keep; // @[BFS.scala 242:21]
  wire  _T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 244:25]
  wire  _select_T_1 = |keep[0]; // @[BFS.scala 250:125]
  wire  _select_T_4 = |keep[1]; // @[BFS.scala 250:125]
  wire  _select_T_7 = |keep[2]; // @[BFS.scala 250:125]
  wire  _select_T_10 = |keep[3]; // @[BFS.scala 250:125]
  wire  _select_T_13 = |keep[4]; // @[BFS.scala 250:125]
  wire  _select_T_16 = |keep[5]; // @[BFS.scala 250:125]
  wire  _select_T_19 = |keep[6]; // @[BFS.scala 250:125]
  wire  _select_T_22 = |keep[7]; // @[BFS.scala 250:125]
  wire  _select_T_25 = |keep[8]; // @[BFS.scala 250:125]
  wire  _select_T_28 = |keep[9]; // @[BFS.scala 250:125]
  wire  _select_T_31 = |keep[10]; // @[BFS.scala 250:125]
  wire  _select_T_34 = |keep[11]; // @[BFS.scala 250:125]
  wire  _select_T_37 = |keep[12]; // @[BFS.scala 250:125]
  wire  _select_T_40 = |keep[13]; // @[BFS.scala 250:125]
  wire  _select_T_43 = |keep[14]; // @[BFS.scala 250:125]
  wire  _select_T_46 = |keep[15]; // @[BFS.scala 250:125]
  wire  _select_T_49 = |keep[16]; // @[BFS.scala 250:125]
  wire  _select_T_52 = |keep[17]; // @[BFS.scala 250:125]
  wire  _select_T_55 = |keep[18]; // @[BFS.scala 250:125]
  wire  _select_T_58 = |keep[19]; // @[BFS.scala 250:125]
  wire  _select_T_61 = |keep[20]; // @[BFS.scala 250:125]
  wire  _select_T_64 = |keep[21]; // @[BFS.scala 250:125]
  wire  _select_T_67 = |keep[22]; // @[BFS.scala 250:125]
  wire  _select_T_70 = |keep[23]; // @[BFS.scala 250:125]
  wire  _select_T_73 = |keep[24]; // @[BFS.scala 250:125]
  wire  _select_T_76 = |keep[25]; // @[BFS.scala 250:125]
  wire  _select_T_79 = |keep[26]; // @[BFS.scala 250:125]
  wire  _select_T_82 = |keep[27]; // @[BFS.scala 250:125]
  wire  _select_T_85 = |keep[28]; // @[BFS.scala 250:125]
  wire  _select_T_88 = |keep[29]; // @[BFS.scala 250:125]
  wire  _select_T_91 = |keep[30]; // @[BFS.scala 250:125]
  wire  _select_T_94 = |keep[31]; // @[BFS.scala 250:125]
  wire [62:0] _select_T_96 = _select_T_94 ? 63'h80000000 : 63'h0; // @[Mux.scala 98:16]
  wire [62:0] _select_T_97 = _select_T_91 ? 63'h40000000 : _select_T_96; // @[Mux.scala 98:16]
  wire [62:0] _select_T_98 = _select_T_88 ? 63'h20000000 : _select_T_97; // @[Mux.scala 98:16]
  wire [62:0] _select_T_99 = _select_T_85 ? 63'h10000000 : _select_T_98; // @[Mux.scala 98:16]
  wire [62:0] _select_T_100 = _select_T_82 ? 63'h8000000 : _select_T_99; // @[Mux.scala 98:16]
  wire [62:0] _select_T_101 = _select_T_79 ? 63'h4000000 : _select_T_100; // @[Mux.scala 98:16]
  wire [62:0] _select_T_102 = _select_T_76 ? 63'h2000000 : _select_T_101; // @[Mux.scala 98:16]
  wire [62:0] _select_T_103 = _select_T_73 ? 63'h1000000 : _select_T_102; // @[Mux.scala 98:16]
  wire [62:0] _select_T_104 = _select_T_70 ? 63'h800000 : _select_T_103; // @[Mux.scala 98:16]
  wire [62:0] _select_T_105 = _select_T_67 ? 63'h400000 : _select_T_104; // @[Mux.scala 98:16]
  wire [62:0] _select_T_106 = _select_T_64 ? 63'h200000 : _select_T_105; // @[Mux.scala 98:16]
  wire [62:0] _select_T_107 = _select_T_61 ? 63'h100000 : _select_T_106; // @[Mux.scala 98:16]
  wire [62:0] _select_T_108 = _select_T_58 ? 63'h80000 : _select_T_107; // @[Mux.scala 98:16]
  wire [62:0] _select_T_109 = _select_T_55 ? 63'h40000 : _select_T_108; // @[Mux.scala 98:16]
  wire [62:0] _select_T_110 = _select_T_52 ? 63'h20000 : _select_T_109; // @[Mux.scala 98:16]
  wire [62:0] _select_T_111 = _select_T_49 ? 63'h10000 : _select_T_110; // @[Mux.scala 98:16]
  wire [62:0] _select_T_112 = _select_T_46 ? 63'h8000 : _select_T_111; // @[Mux.scala 98:16]
  wire [62:0] _select_T_113 = _select_T_43 ? 63'h4000 : _select_T_112; // @[Mux.scala 98:16]
  wire [62:0] _select_T_114 = _select_T_40 ? 63'h2000 : _select_T_113; // @[Mux.scala 98:16]
  wire [62:0] _select_T_115 = _select_T_37 ? 63'h1000 : _select_T_114; // @[Mux.scala 98:16]
  wire [62:0] _select_T_116 = _select_T_34 ? 63'h800 : _select_T_115; // @[Mux.scala 98:16]
  wire [62:0] _select_T_117 = _select_T_31 ? 63'h400 : _select_T_116; // @[Mux.scala 98:16]
  wire [62:0] _select_T_118 = _select_T_28 ? 63'h200 : _select_T_117; // @[Mux.scala 98:16]
  wire [62:0] _select_T_119 = _select_T_25 ? 63'h100 : _select_T_118; // @[Mux.scala 98:16]
  wire [62:0] _select_T_120 = _select_T_22 ? 63'h80 : _select_T_119; // @[Mux.scala 98:16]
  wire [62:0] _select_T_121 = _select_T_19 ? 63'h40 : _select_T_120; // @[Mux.scala 98:16]
  wire [62:0] _select_T_122 = _select_T_16 ? 63'h20 : _select_T_121; // @[Mux.scala 98:16]
  wire [62:0] _select_T_123 = _select_T_13 ? 63'h10 : _select_T_122; // @[Mux.scala 98:16]
  wire [62:0] _select_T_124 = _select_T_10 ? 63'h8 : _select_T_123; // @[Mux.scala 98:16]
  wire [62:0] _select_T_125 = _select_T_7 ? 63'h4 : _select_T_124; // @[Mux.scala 98:16]
  wire [62:0] _select_T_126 = _select_T_4 ? 63'h2 : _select_T_125; // @[Mux.scala 98:16]
  wire [62:0] select = _select_T_1 ? 63'h1 : _select_T_126; // @[Mux.scala 98:16]
  wire [31:0] _io_ddr_out_bits_tdata_T_64 = select[0] ? data[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_65 = select[1] ? data[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_66 = select[2] ? data[95:64] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_67 = select[3] ? data[127:96] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_68 = select[4] ? data[159:128] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_69 = select[5] ? data[191:160] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_70 = select[6] ? data[223:192] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_71 = select[7] ? data[255:224] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_72 = select[8] ? data[287:256] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_73 = select[9] ? data[319:288] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_74 = select[10] ? data[351:320] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_75 = select[11] ? data[383:352] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_76 = select[12] ? data[415:384] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_77 = select[13] ? data[447:416] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_78 = select[14] ? data[479:448] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_79 = select[15] ? data[511:480] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_80 = select[16] ? data[543:512] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_81 = select[17] ? data[575:544] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_82 = select[18] ? data[607:576] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_83 = select[19] ? data[639:608] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_84 = select[20] ? data[671:640] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_85 = select[21] ? data[703:672] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_86 = select[22] ? data[735:704] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_87 = select[23] ? data[767:736] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_88 = select[24] ? data[799:768] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_89 = select[25] ? data[831:800] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_90 = select[26] ? data[863:832] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_91 = select[27] ? data[895:864] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_92 = select[28] ? data[927:896] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_93 = select[29] ? data[959:928] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_94 = select[30] ? data[991:960] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_95 = select[31] ? data[1023:992] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_96 = _io_ddr_out_bits_tdata_T_64 | _io_ddr_out_bits_tdata_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_97 = _io_ddr_out_bits_tdata_T_96 | _io_ddr_out_bits_tdata_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_98 = _io_ddr_out_bits_tdata_T_97 | _io_ddr_out_bits_tdata_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_99 = _io_ddr_out_bits_tdata_T_98 | _io_ddr_out_bits_tdata_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_100 = _io_ddr_out_bits_tdata_T_99 | _io_ddr_out_bits_tdata_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_101 = _io_ddr_out_bits_tdata_T_100 | _io_ddr_out_bits_tdata_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_102 = _io_ddr_out_bits_tdata_T_101 | _io_ddr_out_bits_tdata_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_103 = _io_ddr_out_bits_tdata_T_102 | _io_ddr_out_bits_tdata_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_104 = _io_ddr_out_bits_tdata_T_103 | _io_ddr_out_bits_tdata_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_105 = _io_ddr_out_bits_tdata_T_104 | _io_ddr_out_bits_tdata_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_106 = _io_ddr_out_bits_tdata_T_105 | _io_ddr_out_bits_tdata_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_107 = _io_ddr_out_bits_tdata_T_106 | _io_ddr_out_bits_tdata_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_108 = _io_ddr_out_bits_tdata_T_107 | _io_ddr_out_bits_tdata_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_109 = _io_ddr_out_bits_tdata_T_108 | _io_ddr_out_bits_tdata_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_110 = _io_ddr_out_bits_tdata_T_109 | _io_ddr_out_bits_tdata_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_111 = _io_ddr_out_bits_tdata_T_110 | _io_ddr_out_bits_tdata_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_112 = _io_ddr_out_bits_tdata_T_111 | _io_ddr_out_bits_tdata_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_113 = _io_ddr_out_bits_tdata_T_112 | _io_ddr_out_bits_tdata_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_114 = _io_ddr_out_bits_tdata_T_113 | _io_ddr_out_bits_tdata_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_115 = _io_ddr_out_bits_tdata_T_114 | _io_ddr_out_bits_tdata_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_116 = _io_ddr_out_bits_tdata_T_115 | _io_ddr_out_bits_tdata_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_117 = _io_ddr_out_bits_tdata_T_116 | _io_ddr_out_bits_tdata_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_118 = _io_ddr_out_bits_tdata_T_117 | _io_ddr_out_bits_tdata_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_119 = _io_ddr_out_bits_tdata_T_118 | _io_ddr_out_bits_tdata_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_120 = _io_ddr_out_bits_tdata_T_119 | _io_ddr_out_bits_tdata_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_121 = _io_ddr_out_bits_tdata_T_120 | _io_ddr_out_bits_tdata_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_122 = _io_ddr_out_bits_tdata_T_121 | _io_ddr_out_bits_tdata_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_123 = _io_ddr_out_bits_tdata_T_122 | _io_ddr_out_bits_tdata_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_124 = _io_ddr_out_bits_tdata_T_123 | _io_ddr_out_bits_tdata_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_125 = _io_ddr_out_bits_tdata_T_124 | _io_ddr_out_bits_tdata_T_94; // @[Mux.scala 27:72]
  wire  next_keep_0 = select[0] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_1 = select[1] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_2 = select[2] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_3 = select[3] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_4 = select[4] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_5 = select[5] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_6 = select[6] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_7 = select[7] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_8 = select[8] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_9 = select[9] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_10 = select[10] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_11 = select[11] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_12 = select[12] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_13 = select[13] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_14 = select[14] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_15 = select[15] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_16 = select[16] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_17 = select[17] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_18 = select[18] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_19 = select[19] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_20 = select[20] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_21 = select[21] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_22 = select[22] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_23 = select[23] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_24 = select[24] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_25 = select[25] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_26 = select[26] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_27 = select[27] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_28 = select[28] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_29 = select[29] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_30 = select[30] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_31 = select[31] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire [7:0] keep_lo_lo = {next_keep_7,next_keep_6,next_keep_5,next_keep_4,next_keep_3,next_keep_2,next_keep_1,
    next_keep_0}; // @[BFS.scala 266:36]
  wire [15:0] keep_lo = {next_keep_15,next_keep_14,next_keep_13,next_keep_12,next_keep_11,next_keep_10,next_keep_9,
    next_keep_8,keep_lo_lo}; // @[BFS.scala 266:36]
  wire [7:0] keep_hi_lo = {next_keep_23,next_keep_22,next_keep_21,next_keep_20,next_keep_19,next_keep_18,next_keep_17,
    next_keep_16}; // @[BFS.scala 266:36]
  wire [31:0] _keep_T = {next_keep_31,next_keep_30,next_keep_29,next_keep_28,next_keep_27,next_keep_26,next_keep_25,
    next_keep_24,keep_hi_lo,keep_lo}; // @[BFS.scala 266:36]
  wire [31:0] _keep_T_1 = keep & _keep_T; // @[BFS.scala 266:18]
  assign io_xbar_in_ready = ~(|keep); // @[BFS.scala 247:23]
  assign io_ddr_out_valid = |select; // @[BFS.scala 251:33]
  assign io_ddr_out_bits_tdata = _io_ddr_out_bits_tdata_T_125 | _io_ddr_out_bits_tdata_T_95; // @[Mux.scala 27:72]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 241:21]
      data <= 1024'h0; // @[BFS.scala 241:21]
    end else if (io_xbar_in_valid & io_xbar_in_ready) begin // @[BFS.scala 244:45]
      data <= io_xbar_in_bits_tdata; // @[BFS.scala 245:10]
    end
    if (reset) begin // @[BFS.scala 242:21]
      keep <= 32'h0; // @[BFS.scala 242:21]
    end else if (_T) begin // @[BFS.scala 263:45]
      keep <= io_xbar_in_bits_tkeep; // @[BFS.scala 264:10]
    end else if (io_ddr_out_valid & io_ddr_out_ready) begin // @[BFS.scala 265:52]
      keep <= _keep_T_1; // @[BFS.scala 266:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {32{`RANDOM}};
  data = _RAND_0[1023:0];
  _RAND_1 = {1{`RANDOM}};
  keep = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pipeline_32(
  input         clock,
  input         reset,
  input         io_dout_ready,
  output        io_dout_valid,
  output [31:0] io_dout_bits,
  input         io_din_valid,
  input  [31:0] io_din_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] data; // @[util.scala 238:21]
  reg  valid; // @[util.scala 239:22]
  reg  ready; // @[util.scala 240:22]
  reg [31:0] data2; // @[util.scala 241:22]
  reg  valid2; // @[util.scala 242:23]
  wire  _GEN_1 = ready & io_din_valid; // @[util.scala 247:22 util.scala 249:13 util.scala 252:13]
  assign io_dout_valid = valid; // @[util.scala 268:17]
  assign io_dout_bits = data; // @[util.scala 269:16]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 238:21]
      data <= 32'h0; // @[util.scala 238:21]
    end else if (io_dout_ready) begin // @[util.scala 243:22]
      if (valid2) begin // @[util.scala 244:17]
        data <= data2; // @[util.scala 245:12]
      end else if (ready) begin // @[util.scala 247:22]
        data <= io_din_bits; // @[util.scala 248:12]
      end else begin
        data <= 32'h0; // @[util.scala 251:12]
      end
    end
    if (reset) begin // @[util.scala 239:22]
      valid <= 1'h0; // @[util.scala 239:22]
    end else if (io_dout_ready) begin // @[util.scala 243:22]
      if (valid2) begin // @[util.scala 244:17]
        valid <= valid2; // @[util.scala 246:13]
      end else begin
        valid <= _GEN_1;
      end
    end
    if (reset) begin // @[util.scala 240:22]
      ready <= 1'h0; // @[util.scala 240:22]
    end else begin
      ready <= io_dout_ready; // @[util.scala 255:9]
    end
    if (reset) begin // @[util.scala 241:22]
      data2 <= 32'h0; // @[util.scala 241:22]
    end else if (~io_dout_ready & ready) begin // @[util.scala 258:33]
      data2 <= io_din_bits; // @[util.scala 259:11]
    end else if (io_dout_ready) begin // @[util.scala 261:28]
      data2 <= 32'h0; // @[util.scala 263:11]
    end
    if (reset) begin // @[util.scala 242:23]
      valid2 <= 1'h0; // @[util.scala 242:23]
    end else if (~io_dout_ready & ready) begin // @[util.scala 258:33]
      valid2 <= io_din_valid; // @[util.scala 260:12]
    end else if (io_dout_ready) begin // @[util.scala 261:28]
      valid2 <= 1'h0; // @[util.scala 264:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ready = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  data2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  valid2 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pipeline_34(
  input        clock,
  input        reset,
  input        io_dout_ready,
  output       io_dout_valid,
  output [8:0] io_dout_bits,
  input        io_din_valid,
  input  [8:0] io_din_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] data; // @[util.scala 238:21]
  reg  valid; // @[util.scala 239:22]
  reg  ready; // @[util.scala 240:22]
  reg [8:0] data2; // @[util.scala 241:22]
  reg  valid2; // @[util.scala 242:23]
  wire  _GEN_1 = ready & io_din_valid; // @[util.scala 247:22 util.scala 249:13 util.scala 252:13]
  assign io_dout_valid = valid; // @[util.scala 268:17]
  assign io_dout_bits = data; // @[util.scala 269:16]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 238:21]
      data <= 9'h0; // @[util.scala 238:21]
    end else if (io_dout_ready) begin // @[util.scala 243:22]
      if (valid2) begin // @[util.scala 244:17]
        data <= data2; // @[util.scala 245:12]
      end else if (ready) begin // @[util.scala 247:22]
        data <= io_din_bits; // @[util.scala 248:12]
      end else begin
        data <= 9'h0; // @[util.scala 251:12]
      end
    end
    if (reset) begin // @[util.scala 239:22]
      valid <= 1'h0; // @[util.scala 239:22]
    end else if (io_dout_ready) begin // @[util.scala 243:22]
      if (valid2) begin // @[util.scala 244:17]
        valid <= valid2; // @[util.scala 246:13]
      end else begin
        valid <= _GEN_1;
      end
    end
    if (reset) begin // @[util.scala 240:22]
      ready <= 1'h0; // @[util.scala 240:22]
    end else begin
      ready <= io_dout_ready; // @[util.scala 255:9]
    end
    if (reset) begin // @[util.scala 241:22]
      data2 <= 9'h0; // @[util.scala 241:22]
    end else if (~io_dout_ready & ready) begin // @[util.scala 258:33]
      data2 <= io_din_bits; // @[util.scala 259:11]
    end else if (io_dout_ready) begin // @[util.scala 261:28]
      data2 <= 9'h0; // @[util.scala 263:11]
    end
    if (reset) begin // @[util.scala 242:23]
      valid2 <= 1'h0; // @[util.scala 242:23]
    end else if (~io_dout_ready & ready) begin // @[util.scala 258:33]
      valid2 <= io_din_valid; // @[util.scala 260:12]
    end else if (io_dout_ready) begin // @[util.scala 261:28]
      valid2 <= 1'h0; // @[util.scala 264:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ready = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  data2 = _RAND_3[8:0];
  _RAND_4 = {1{`RANDOM}};
  valid2 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Scatter(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h0 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h0 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h0 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h0 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h0 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h0 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h0 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h0 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h0 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h0 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h0 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h0 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h0 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h0 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h0 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h0 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h0 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h0 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h0 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h0 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h0 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h0 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h0 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h0 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h0 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h0 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h0 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h0 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h0 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h0 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h0 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h0 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_1(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h1 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h1 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h1 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h1 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h1 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h1 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h1 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h1 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h1 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h1 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h1 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h1 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h1 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h1 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h1 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h1 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h1 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h1 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h1 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h1 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h1 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h1 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h1 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h1 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h1 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h1 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h1 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h1 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h1 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h1 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h1 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h1 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_2(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h2 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h2 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h2 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h2 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h2 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h2 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h2 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h2 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h2 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h2 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h2 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h2 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h2 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h2 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h2 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h2 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h2 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h2 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h2 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h2 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h2 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h2 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h2 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h2 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h2 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h2 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h2 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h2 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h2 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h2 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h2 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h2 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_3(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h3 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h3 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h3 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h3 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h3 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h3 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h3 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h3 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h3 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h3 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h3 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h3 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h3 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h3 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h3 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h3 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h3 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h3 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h3 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h3 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h3 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h3 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h3 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h3 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h3 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h3 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h3 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h3 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h3 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h3 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h3 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h3 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_4(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h4 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h4 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h4 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h4 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h4 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h4 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h4 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h4 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h4 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h4 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h4 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h4 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h4 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h4 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h4 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h4 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h4 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h4 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h4 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h4 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h4 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h4 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h4 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h4 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h4 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h4 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h4 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h4 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h4 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h4 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h4 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h4 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_5(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h5 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h5 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h5 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h5 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h5 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h5 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h5 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h5 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h5 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h5 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h5 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h5 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h5 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h5 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h5 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h5 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h5 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h5 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h5 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h5 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h5 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h5 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h5 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h5 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h5 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h5 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h5 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h5 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h5 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h5 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h5 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h5 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_6(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h6 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h6 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h6 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h6 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h6 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h6 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h6 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h6 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h6 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h6 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h6 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h6 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h6 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h6 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h6 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h6 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h6 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h6 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h6 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h6 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h6 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h6 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h6 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h6 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h6 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h6 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h6 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h6 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h6 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h6 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h6 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h6 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_7(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h7 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h7 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h7 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h7 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h7 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h7 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h7 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h7 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h7 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h7 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h7 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h7 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h7 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h7 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h7 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h7 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h7 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h7 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h7 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h7 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h7 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h7 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h7 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h7 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h7 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h7 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h7 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h7 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h7 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h7 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h7 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h7 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_8(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h8 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h8 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h8 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h8 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h8 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h8 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h8 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h8 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h8 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h8 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h8 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h8 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h8 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h8 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h8 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h8 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h8 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h8 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h8 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h8 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h8 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h8 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h8 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h8 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h8 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h8 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h8 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h8 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h8 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h8 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h8 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h8 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_9(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'h9 & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'h9 & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'h9 & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'h9 & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'h9 & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'h9 & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'h9 & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'h9 & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'h9 & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'h9 & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'h9 & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'h9 & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'h9 & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'h9 & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'h9 & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'h9 & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'h9 & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'h9 & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'h9 & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'h9 & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'h9 & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'h9 & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'h9 & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'h9 & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'h9 & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'h9 & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'h9 & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'h9 & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'h9 & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'h9 & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'h9 & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'h9 & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_10(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'ha & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'ha & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'ha & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'ha & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'ha & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'ha & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'ha & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'ha & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'ha & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'ha & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'ha & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'ha & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'ha & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'ha & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'ha & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'ha & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'ha & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'ha & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'ha & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'ha & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'ha & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'ha & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'ha & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'ha & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'ha & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'ha & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'ha & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'ha & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'ha & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'ha & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'ha & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'ha & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_11(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'hb & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'hb & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'hb & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'hb & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'hb & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'hb & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'hb & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'hb & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'hb & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'hb & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'hb & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'hb & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'hb & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'hb & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'hb & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'hb & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'hb & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'hb & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'hb & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'hb & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'hb & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'hb & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'hb & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'hb & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'hb & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'hb & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'hb & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'hb & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'hb & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'hb & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'hb & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'hb & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_12(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'hc & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'hc & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'hc & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'hc & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'hc & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'hc & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'hc & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'hc & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'hc & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'hc & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'hc & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'hc & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'hc & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'hc & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'hc & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'hc & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'hc & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'hc & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'hc & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'hc & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'hc & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'hc & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'hc & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'hc & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'hc & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'hc & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'hc & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'hc & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'hc & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'hc & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'hc & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'hc & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_13(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'hd & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'hd & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'hd & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'hd & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'hd & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'hd & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'hd & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'hd & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'hd & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'hd & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'hd & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'hd & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'hd & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'hd & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'hd & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'hd & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'hd & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'hd & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'hd & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'hd & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'hd & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'hd & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'hd & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'hd & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'hd & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'hd & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'hd & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'hd & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'hd & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'hd & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'hd & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'hd & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_14(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'he & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'he & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'he & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'he & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'he & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'he & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'he & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'he & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'he & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'he & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'he & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'he & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'he & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'he & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'he & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'he & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'he & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'he & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'he & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'he & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'he & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'he & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'he & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'he & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'he & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'he & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'he & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'he & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'he & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'he & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'he & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'he & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module Scatter_15(
  input           clock,
  input           reset,
  output          io_xbar_in_ready,
  input           io_xbar_in_valid,
  input  [1023:0] io_xbar_in_bits_tdata,
  input  [31:0]   io_xbar_in_bits_tkeep,
  input           io_ddr_out_ready,
  output          io_ddr_out_valid,
  output [31:0]   io_ddr_out_bits_tdata,
  output          io_end,
  input           io_local_fpga_id
);
  wire [16:0] bitmap__addra; // @[BFS.scala 699:22]
  wire  bitmap__clka; // @[BFS.scala 699:22]
  wire [8:0] bitmap__dina; // @[BFS.scala 699:22]
  wire  bitmap__ena; // @[BFS.scala 699:22]
  wire  bitmap__wea; // @[BFS.scala 699:22]
  wire [16:0] bitmap__addrb; // @[BFS.scala 699:22]
  wire  bitmap__clkb; // @[BFS.scala 699:22]
  wire [8:0] bitmap__doutb; // @[BFS.scala 699:22]
  wire  bitmap__enb; // @[BFS.scala 699:22]
  wire  arbi_clock; // @[BFS.scala 700:20]
  wire  arbi_reset; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_ready; // @[BFS.scala 700:20]
  wire  arbi_io_xbar_in_valid; // @[BFS.scala 700:20]
  wire [1023:0] arbi_io_xbar_in_bits_tdata; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_xbar_in_bits_tkeep; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_ready; // @[BFS.scala 700:20]
  wire  arbi_io_ddr_out_valid; // @[BFS.scala 700:20]
  wire [31:0] arbi_io_ddr_out_bits_tdata; // @[BFS.scala 700:20]
  wire  vertex_in_fifo_full; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_din; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_wr_en; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_empty; // @[BFS.scala 738:30]
  wire [31:0] vertex_in_fifo_dout; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_rd_en; // @[BFS.scala 738:30]
  wire [5:0] vertex_in_fifo_data_count; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_clk; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_srst; // @[BFS.scala 738:30]
  wire  vertex_in_fifo_valid; // @[BFS.scala 738:30]
  wire  vertex_out_fifo_full; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_din; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 739:31]
  wire [31:0] vertex_out_fifo_dout; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 739:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 739:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 739:31]
  wire  bitmap_wait_clock; // @[BFS.scala 748:27]
  wire  bitmap_wait_reset; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_ready; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_dout_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_dout_bits; // @[BFS.scala 748:27]
  wire  bitmap_wait_io_din_valid; // @[BFS.scala 748:27]
  wire [31:0] bitmap_wait_io_din_bits; // @[BFS.scala 748:27]
  wire  bitmap_write_addr_clock; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_reset; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_ready; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_dout_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_dout_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_addr_io_din_valid; // @[BFS.scala 753:33]
  wire [31:0] bitmap_write_addr_io_din_bits; // @[BFS.scala 753:33]
  wire  bitmap_write_data_clock; // @[BFS.scala 758:33]
  wire  bitmap_write_data_reset; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_ready; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_dout_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_dout_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_io_din_valid; // @[BFS.scala 758:33]
  wire [8:0] bitmap_write_data_io_din_bits; // @[BFS.scala 758:33]
  wire  bitmap_write_data_forward_clock; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_reset; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_ready; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_dout_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_dout_bits; // @[BFS.scala 763:41]
  wire  bitmap_write_data_forward_io_din_valid; // @[BFS.scala 763:41]
  wire [8:0] bitmap_write_data_forward_io_din_bits; // @[BFS.scala 763:41]
  wire  _filtered_keep_0_T_7 = io_xbar_in_bits_tdata[4] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_0_T_8 = io_xbar_in_bits_tdata[3:0] == 4'hf & _filtered_keep_0_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_0_T_9 = io_xbar_in_bits_tdata[31] | _filtered_keep_0_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_1_T_7 = io_xbar_in_bits_tdata[36] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_1_T_8 = io_xbar_in_bits_tdata[35:32] == 4'hf & _filtered_keep_1_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_1_T_9 = io_xbar_in_bits_tdata[63] | _filtered_keep_1_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_2_T_7 = io_xbar_in_bits_tdata[68] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_2_T_8 = io_xbar_in_bits_tdata[67:64] == 4'hf & _filtered_keep_2_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_2_T_9 = io_xbar_in_bits_tdata[95] | _filtered_keep_2_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_3_T_7 = io_xbar_in_bits_tdata[100] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_3_T_8 = io_xbar_in_bits_tdata[99:96] == 4'hf & _filtered_keep_3_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_3_T_9 = io_xbar_in_bits_tdata[127] | _filtered_keep_3_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_4_T_7 = io_xbar_in_bits_tdata[132] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_4_T_8 = io_xbar_in_bits_tdata[131:128] == 4'hf & _filtered_keep_4_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_4_T_9 = io_xbar_in_bits_tdata[159] | _filtered_keep_4_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_5_T_7 = io_xbar_in_bits_tdata[164] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_5_T_8 = io_xbar_in_bits_tdata[163:160] == 4'hf & _filtered_keep_5_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_5_T_9 = io_xbar_in_bits_tdata[191] | _filtered_keep_5_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_6_T_7 = io_xbar_in_bits_tdata[196] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_6_T_8 = io_xbar_in_bits_tdata[195:192] == 4'hf & _filtered_keep_6_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_6_T_9 = io_xbar_in_bits_tdata[223] | _filtered_keep_6_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_7_T_7 = io_xbar_in_bits_tdata[228] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_7_T_8 = io_xbar_in_bits_tdata[227:224] == 4'hf & _filtered_keep_7_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_7_T_9 = io_xbar_in_bits_tdata[255] | _filtered_keep_7_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_8_T_7 = io_xbar_in_bits_tdata[260] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_8_T_8 = io_xbar_in_bits_tdata[259:256] == 4'hf & _filtered_keep_8_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_8_T_9 = io_xbar_in_bits_tdata[287] | _filtered_keep_8_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_9_T_7 = io_xbar_in_bits_tdata[292] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_9_T_8 = io_xbar_in_bits_tdata[291:288] == 4'hf & _filtered_keep_9_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_9_T_9 = io_xbar_in_bits_tdata[319] | _filtered_keep_9_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_10_T_7 = io_xbar_in_bits_tdata[324] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_10_T_8 = io_xbar_in_bits_tdata[323:320] == 4'hf & _filtered_keep_10_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_10_T_9 = io_xbar_in_bits_tdata[351] | _filtered_keep_10_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_11_T_7 = io_xbar_in_bits_tdata[356] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_11_T_8 = io_xbar_in_bits_tdata[355:352] == 4'hf & _filtered_keep_11_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_11_T_9 = io_xbar_in_bits_tdata[383] | _filtered_keep_11_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_12_T_7 = io_xbar_in_bits_tdata[388] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_12_T_8 = io_xbar_in_bits_tdata[387:384] == 4'hf & _filtered_keep_12_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_12_T_9 = io_xbar_in_bits_tdata[415] | _filtered_keep_12_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_13_T_7 = io_xbar_in_bits_tdata[420] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_13_T_8 = io_xbar_in_bits_tdata[419:416] == 4'hf & _filtered_keep_13_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_13_T_9 = io_xbar_in_bits_tdata[447] | _filtered_keep_13_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_14_T_7 = io_xbar_in_bits_tdata[452] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_14_T_8 = io_xbar_in_bits_tdata[451:448] == 4'hf & _filtered_keep_14_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_14_T_9 = io_xbar_in_bits_tdata[479] | _filtered_keep_14_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_15_T_7 = io_xbar_in_bits_tdata[484] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_15_T_8 = io_xbar_in_bits_tdata[483:480] == 4'hf & _filtered_keep_15_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_15_T_9 = io_xbar_in_bits_tdata[511] | _filtered_keep_15_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_16_T_7 = io_xbar_in_bits_tdata[516] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_16_T_8 = io_xbar_in_bits_tdata[515:512] == 4'hf & _filtered_keep_16_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_16_T_9 = io_xbar_in_bits_tdata[543] | _filtered_keep_16_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_16 = io_xbar_in_bits_tkeep[16] & _filtered_keep_16_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_17_T_7 = io_xbar_in_bits_tdata[548] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_17_T_8 = io_xbar_in_bits_tdata[547:544] == 4'hf & _filtered_keep_17_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_17_T_9 = io_xbar_in_bits_tdata[575] | _filtered_keep_17_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_17 = io_xbar_in_bits_tkeep[17] & _filtered_keep_17_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_18_T_7 = io_xbar_in_bits_tdata[580] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_18_T_8 = io_xbar_in_bits_tdata[579:576] == 4'hf & _filtered_keep_18_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_18_T_9 = io_xbar_in_bits_tdata[607] | _filtered_keep_18_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_18 = io_xbar_in_bits_tkeep[18] & _filtered_keep_18_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_19_T_7 = io_xbar_in_bits_tdata[612] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_19_T_8 = io_xbar_in_bits_tdata[611:608] == 4'hf & _filtered_keep_19_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_19_T_9 = io_xbar_in_bits_tdata[639] | _filtered_keep_19_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_19 = io_xbar_in_bits_tkeep[19] & _filtered_keep_19_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_20_T_7 = io_xbar_in_bits_tdata[644] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_20_T_8 = io_xbar_in_bits_tdata[643:640] == 4'hf & _filtered_keep_20_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_20_T_9 = io_xbar_in_bits_tdata[671] | _filtered_keep_20_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_20 = io_xbar_in_bits_tkeep[20] & _filtered_keep_20_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_21_T_7 = io_xbar_in_bits_tdata[676] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_21_T_8 = io_xbar_in_bits_tdata[675:672] == 4'hf & _filtered_keep_21_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_21_T_9 = io_xbar_in_bits_tdata[703] | _filtered_keep_21_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_21 = io_xbar_in_bits_tkeep[21] & _filtered_keep_21_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_22_T_7 = io_xbar_in_bits_tdata[708] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_22_T_8 = io_xbar_in_bits_tdata[707:704] == 4'hf & _filtered_keep_22_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_22_T_9 = io_xbar_in_bits_tdata[735] | _filtered_keep_22_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_22 = io_xbar_in_bits_tkeep[22] & _filtered_keep_22_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_23_T_7 = io_xbar_in_bits_tdata[740] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_23_T_8 = io_xbar_in_bits_tdata[739:736] == 4'hf & _filtered_keep_23_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_23_T_9 = io_xbar_in_bits_tdata[767] | _filtered_keep_23_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_23 = io_xbar_in_bits_tkeep[23] & _filtered_keep_23_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_24_T_7 = io_xbar_in_bits_tdata[772] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_24_T_8 = io_xbar_in_bits_tdata[771:768] == 4'hf & _filtered_keep_24_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_24_T_9 = io_xbar_in_bits_tdata[799] | _filtered_keep_24_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_24 = io_xbar_in_bits_tkeep[24] & _filtered_keep_24_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_25_T_7 = io_xbar_in_bits_tdata[804] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_25_T_8 = io_xbar_in_bits_tdata[803:800] == 4'hf & _filtered_keep_25_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_25_T_9 = io_xbar_in_bits_tdata[831] | _filtered_keep_25_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_25 = io_xbar_in_bits_tkeep[25] & _filtered_keep_25_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_26_T_7 = io_xbar_in_bits_tdata[836] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_26_T_8 = io_xbar_in_bits_tdata[835:832] == 4'hf & _filtered_keep_26_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_26_T_9 = io_xbar_in_bits_tdata[863] | _filtered_keep_26_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_26 = io_xbar_in_bits_tkeep[26] & _filtered_keep_26_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_27_T_7 = io_xbar_in_bits_tdata[868] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_27_T_8 = io_xbar_in_bits_tdata[867:864] == 4'hf & _filtered_keep_27_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_27_T_9 = io_xbar_in_bits_tdata[895] | _filtered_keep_27_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_27 = io_xbar_in_bits_tkeep[27] & _filtered_keep_27_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_28_T_7 = io_xbar_in_bits_tdata[900] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_28_T_8 = io_xbar_in_bits_tdata[899:896] == 4'hf & _filtered_keep_28_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_28_T_9 = io_xbar_in_bits_tdata[927] | _filtered_keep_28_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_28 = io_xbar_in_bits_tkeep[28] & _filtered_keep_28_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_29_T_7 = io_xbar_in_bits_tdata[932] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_29_T_8 = io_xbar_in_bits_tdata[931:928] == 4'hf & _filtered_keep_29_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_29_T_9 = io_xbar_in_bits_tdata[959] | _filtered_keep_29_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_29 = io_xbar_in_bits_tkeep[29] & _filtered_keep_29_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_30_T_7 = io_xbar_in_bits_tdata[964] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_30_T_8 = io_xbar_in_bits_tdata[963:960] == 4'hf & _filtered_keep_30_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_30_T_9 = io_xbar_in_bits_tdata[991] | _filtered_keep_30_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_30 = io_xbar_in_bits_tkeep[30] & _filtered_keep_30_T_9; // @[BFS.scala 726:15]
  wire  _filtered_keep_31_T_7 = io_xbar_in_bits_tdata[996] == io_local_fpga_id; // @[BFS.scala 707:80]
  wire  _filtered_keep_31_T_8 = io_xbar_in_bits_tdata[995:992] == 4'hf & _filtered_keep_31_T_7; // @[BFS.scala 706:47]
  wire  _filtered_keep_31_T_9 = io_xbar_in_bits_tdata[1023] | _filtered_keep_31_T_8; // @[BFS.scala 727:12]
  wire  filtered_keep_31 = io_xbar_in_bits_tkeep[31] & _filtered_keep_31_T_9; // @[BFS.scala 726:15]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_lo_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_lo = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,arbi_io_xbar_in_bits_tkeep_lo_lo}; // @[BFS.scala 732:53]
  wire [7:0] arbi_io_xbar_in_bits_tkeep_hi_lo = {filtered_keep_23,filtered_keep_22,filtered_keep_21,filtered_keep_20,
    filtered_keep_19,filtered_keep_18,filtered_keep_17,filtered_keep_16}; // @[BFS.scala 732:53]
  wire [15:0] arbi_io_xbar_in_bits_tkeep_hi = {filtered_keep_31,filtered_keep_30,filtered_keep_29,filtered_keep_28,
    filtered_keep_27,filtered_keep_26,filtered_keep_25,filtered_keep_24,arbi_io_xbar_in_bits_tkeep_hi_lo}; // @[BFS.scala 732:53]
  wire  halt = vertex_out_fifo_full; // @[BFS.scala 747:38]
  wire [26:0] _GEN_0 = {{1'd0}, bitmap_wait_io_dout_bits[30:5]}; // @[BFS.scala 718:59]
  wire  _bitmap_write_addr_io_din_valid_T_1 = _GEN_0 > 27'he7fff; // @[BFS.scala 718:59]
  wire [3:0] _bitmap_write_addr_io_din_valid_WIRE = {{1'd0}, bitmap_wait_io_dout_bits[7:5]}; // @[BFS.scala 720:107 BFS.scala 720:107]
  wire [3:0] _bitmap_write_addr_io_din_valid_T_3 = _GEN_0 > 27'he7fff ? 4'h8 : _bitmap_write_addr_io_din_valid_WIRE; // @[BFS.scala 718:8]
  wire [26:0] _bitmap_doutb_T_5 = _GEN_0 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE = {{4'd0}, bitmap_wait_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_7 = _bitmap_write_addr_io_din_valid_T_1 ? _bitmap_doutb_T_5 : _bitmap_doutb_WIRE; // @[BFS.scala 712:8]
  wire [26:0] _GEN_3 = {{1'd0}, bitmap_write_addr_io_dout_bits[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_doutb_T_12 = _GEN_3 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_doutb_WIRE_1 = {{4'd0}, bitmap_write_addr_io_dout_bits[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_doutb_T_14 = _GEN_3 > 27'he7fff ? _bitmap_doutb_T_12 : _bitmap_doutb_WIRE_1; // @[BFS.scala 712:8]
  wire  _bitmap_doutb_T_15 = _bitmap_doutb_T_7 == _bitmap_doutb_T_14; // @[BFS.scala 770:49]
  wire  _bitmap_doutb_T_16 = bitmap_write_addr_io_dout_valid & bitmap_wait_io_dout_valid & _bitmap_doutb_T_15; // @[BFS.scala 769:67]
  wire [8:0] _bitmap_doutb_T_17 = bitmap_write_data_forward_io_dout_valid ? bitmap_write_data_forward_io_dout_bits :
    bitmap__doutb; // @[Mux.scala 98:16]
  wire [8:0] bitmap_doutb = _bitmap_doutb_T_16 ? bitmap_write_data_io_dout_bits : _bitmap_doutb_T_17; // @[Mux.scala 98:16]
  wire [8:0] _bitmap_write_addr_io_din_valid_T_4 = bitmap_doutb >> _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 755:18]
  wire  _bitmap_write_addr_io_din_valid_T_9 = ~_bitmap_write_addr_io_din_valid_T_4[0] | bitmap_wait_io_dout_bits[31]; // @[BFS.scala 755:77]
  wire [23:0] _bitmap_write_data_io_din_bits_T_4 = 24'h1 << _bitmap_write_addr_io_din_valid_T_3; // @[BFS.scala 761:61]
  wire [23:0] _GEN_7 = {{15'd0}, bitmap_doutb}; // @[BFS.scala 761:49]
  wire [23:0] _bitmap_write_data_io_din_bits_T_5 = _GEN_7 | _bitmap_write_data_io_din_bits_T_4; // @[BFS.scala 761:49]
  wire [26:0] _GEN_8 = {{1'd0}, vertex_in_fifo_dout[30:5]}; // @[BFS.scala 712:59]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_5 = _GEN_8 - 27'he7fff; // @[BFS.scala 713:57]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_WIRE = {{4'd0}, vertex_in_fifo_dout[30:8]}; // @[BFS.scala 714:69 BFS.scala 714:69]
  wire [26:0] _bitmap_write_data_forward_io_din_valid_T_7 = _GEN_8 > 27'he7fff ?
    _bitmap_write_data_forward_io_din_valid_T_5 : _bitmap_write_data_forward_io_din_valid_WIRE; // @[BFS.scala 712:8]
  wire  _bitmap_write_data_forward_io_din_valid_T_15 = _bitmap_write_data_forward_io_din_valid_T_7 == _bitmap_doutb_T_14
    ; // @[BFS.scala 765:46]
  wire [31:0] _io_end_T = {{31'd0}, vertex_out_fifo_dout[31]}; // @[util.scala 207:12]
  bitmap_0 bitmap_ ( // @[BFS.scala 699:22]
    .addra(bitmap__addra),
    .clka(bitmap__clka),
    .dina(bitmap__dina),
    .ena(bitmap__ena),
    .wea(bitmap__wea),
    .addrb(bitmap__addrb),
    .clkb(bitmap__clkb),
    .doutb(bitmap__doutb),
    .enb(bitmap__enb)
  );
  axis_arbitrator arbi ( // @[BFS.scala 700:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_xbar_in_ready(arbi_io_xbar_in_ready),
    .io_xbar_in_valid(arbi_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(arbi_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(arbi_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(arbi_io_ddr_out_ready),
    .io_ddr_out_valid(arbi_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(arbi_io_ddr_out_bits_tdata)
  );
  vid_fifo vertex_in_fifo ( // @[BFS.scala 738:30]
    .full(vertex_in_fifo_full),
    .din(vertex_in_fifo_din),
    .wr_en(vertex_in_fifo_wr_en),
    .empty(vertex_in_fifo_empty),
    .dout(vertex_in_fifo_dout),
    .rd_en(vertex_in_fifo_rd_en),
    .data_count(vertex_in_fifo_data_count),
    .clk(vertex_in_fifo_clk),
    .srst(vertex_in_fifo_srst),
    .valid(vertex_in_fifo_valid)
  );
  vid_fifo vertex_out_fifo ( // @[BFS.scala 739:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  pipeline_32 bitmap_wait ( // @[BFS.scala 748:27]
    .clock(bitmap_wait_clock),
    .reset(bitmap_wait_reset),
    .io_dout_ready(bitmap_wait_io_dout_ready),
    .io_dout_valid(bitmap_wait_io_dout_valid),
    .io_dout_bits(bitmap_wait_io_dout_bits),
    .io_din_valid(bitmap_wait_io_din_valid),
    .io_din_bits(bitmap_wait_io_din_bits)
  );
  pipeline_32 bitmap_write_addr ( // @[BFS.scala 753:33]
    .clock(bitmap_write_addr_clock),
    .reset(bitmap_write_addr_reset),
    .io_dout_ready(bitmap_write_addr_io_dout_ready),
    .io_dout_valid(bitmap_write_addr_io_dout_valid),
    .io_dout_bits(bitmap_write_addr_io_dout_bits),
    .io_din_valid(bitmap_write_addr_io_din_valid),
    .io_din_bits(bitmap_write_addr_io_din_bits)
  );
  pipeline_34 bitmap_write_data ( // @[BFS.scala 758:33]
    .clock(bitmap_write_data_clock),
    .reset(bitmap_write_data_reset),
    .io_dout_ready(bitmap_write_data_io_dout_ready),
    .io_dout_valid(bitmap_write_data_io_dout_valid),
    .io_dout_bits(bitmap_write_data_io_dout_bits),
    .io_din_valid(bitmap_write_data_io_din_valid),
    .io_din_bits(bitmap_write_data_io_din_bits)
  );
  pipeline_34 bitmap_write_data_forward ( // @[BFS.scala 763:41]
    .clock(bitmap_write_data_forward_clock),
    .reset(bitmap_write_data_forward_reset),
    .io_dout_ready(bitmap_write_data_forward_io_dout_ready),
    .io_dout_valid(bitmap_write_data_forward_io_dout_valid),
    .io_dout_bits(bitmap_write_data_forward_io_dout_bits),
    .io_din_valid(bitmap_write_data_forward_io_din_valid),
    .io_din_bits(bitmap_write_data_forward_io_din_bits)
  );
  assign io_xbar_in_ready = arbi_io_xbar_in_ready; // @[BFS.scala 736:20]
  assign io_ddr_out_valid = vertex_out_fifo_valid & ~vertex_out_fifo_dout[31]; // @[BFS.scala 789:50]
  assign io_ddr_out_bits_tdata = vertex_out_fifo_dout; // @[BFS.scala 792:25]
  assign io_end = _io_end_T[0] & ~vertex_out_fifo_empty; // @[util.scala 207:36]
  assign bitmap__addra = _bitmap_doutb_T_14[16:0]; // @[BFS.scala 787:19]
  assign bitmap__clka = clock; // @[BFS.scala 785:33]
  assign bitmap__dina = bitmap_write_data_io_dout_bits; // @[BFS.scala 786:18]
  assign bitmap__ena = 1'h1; // @[BFS.scala 783:17]
  assign bitmap__wea = bitmap_write_addr_io_dout_valid & ~bitmap_write_addr_io_dout_bits[31]; // @[BFS.scala 784:52]
  assign bitmap__addrb = _bitmap_write_data_forward_io_din_valid_T_7[16:0]; // @[BFS.scala 778:19]
  assign bitmap__clkb = clock; // @[BFS.scala 779:33]
  assign bitmap__enb = 1'h1; // @[BFS.scala 777:17]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_xbar_in_valid = io_xbar_in_valid; // @[BFS.scala 734:25]
  assign arbi_io_xbar_in_bits_tdata = io_xbar_in_bits_tdata; // @[BFS.scala 733:30]
  assign arbi_io_xbar_in_bits_tkeep = {arbi_io_xbar_in_bits_tkeep_hi,arbi_io_xbar_in_bits_tkeep_lo}; // @[BFS.scala 732:53]
  assign arbi_io_ddr_out_ready = ~vertex_in_fifo_full; // @[BFS.scala 776:51]
  assign vertex_in_fifo_din = arbi_io_ddr_out_bits_tdata; // @[BFS.scala 774:25]
  assign vertex_in_fifo_wr_en = arbi_io_ddr_out_valid; // @[BFS.scala 775:27]
  assign vertex_in_fifo_rd_en = ~halt; // @[BFS.scala 780:30]
  assign vertex_in_fifo_clk = clock; // @[BFS.scala 740:40]
  assign vertex_in_fifo_srst = reset; // @[BFS.scala 741:41]
  assign vertex_out_fifo_din = bitmap_write_addr_io_dout_bits; // @[BFS.scala 782:26]
  assign vertex_out_fifo_wr_en = bitmap_write_addr_io_dout_valid; // @[BFS.scala 781:28]
  assign vertex_out_fifo_rd_en = io_ddr_out_ready; // @[BFS.scala 788:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 742:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 743:42]
  assign bitmap_wait_clock = clock;
  assign bitmap_wait_reset = reset;
  assign bitmap_wait_io_dout_ready = ~halt; // @[BFS.scala 751:32]
  assign bitmap_wait_io_din_valid = vertex_in_fifo_valid; // @[BFS.scala 749:28]
  assign bitmap_wait_io_din_bits = vertex_in_fifo_dout; // @[BFS.scala 750:27]
  assign bitmap_write_addr_clock = clock;
  assign bitmap_write_addr_reset = reset;
  assign bitmap_write_addr_io_dout_ready = ~halt; // @[BFS.scala 757:38]
  assign bitmap_write_addr_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 754:63]
  assign bitmap_write_addr_io_din_bits = bitmap_wait_io_dout_bits; // @[BFS.scala 756:33]
  assign bitmap_write_data_clock = clock;
  assign bitmap_write_data_reset = reset;
  assign bitmap_write_data_io_dout_ready = ~halt; // @[BFS.scala 762:38]
  assign bitmap_write_data_io_din_valid = bitmap_wait_io_dout_valid & _bitmap_write_addr_io_din_valid_T_9; // @[BFS.scala 759:64]
  assign bitmap_write_data_io_din_bits = _bitmap_write_data_io_din_bits_T_5[8:0]; // @[BFS.scala 761:33]
  assign bitmap_write_data_forward_clock = clock;
  assign bitmap_write_data_forward_reset = reset;
  assign bitmap_write_data_forward_io_dout_ready = ~halt; // @[BFS.scala 767:46]
  assign bitmap_write_data_forward_io_din_valid = bitmap_write_addr_io_dout_valid & vertex_in_fifo_valid &
    _bitmap_write_data_forward_io_din_valid_T_15; // @[BFS.scala 764:95]
  assign bitmap_write_data_forward_io_din_bits = bitmap_write_data_io_dout_bits; // @[BFS.scala 766:41]
endmodule
module axis_arbitrator_16(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] data; // @[BFS.scala 241:21]
  reg [15:0] keep; // @[BFS.scala 242:21]
  wire  _T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 244:25]
  wire  _select_T_1 = |keep[0]; // @[BFS.scala 250:125]
  wire  _select_T_4 = |keep[1]; // @[BFS.scala 250:125]
  wire  _select_T_7 = |keep[2]; // @[BFS.scala 250:125]
  wire  _select_T_10 = |keep[3]; // @[BFS.scala 250:125]
  wire  _select_T_13 = |keep[4]; // @[BFS.scala 250:125]
  wire  _select_T_16 = |keep[5]; // @[BFS.scala 250:125]
  wire  _select_T_19 = |keep[6]; // @[BFS.scala 250:125]
  wire  _select_T_22 = |keep[7]; // @[BFS.scala 250:125]
  wire  _select_T_25 = |keep[8]; // @[BFS.scala 250:125]
  wire  _select_T_28 = |keep[9]; // @[BFS.scala 250:125]
  wire  _select_T_31 = |keep[10]; // @[BFS.scala 250:125]
  wire  _select_T_34 = |keep[11]; // @[BFS.scala 250:125]
  wire  _select_T_37 = |keep[12]; // @[BFS.scala 250:125]
  wire  _select_T_40 = |keep[13]; // @[BFS.scala 250:125]
  wire  _select_T_43 = |keep[14]; // @[BFS.scala 250:125]
  wire  _select_T_46 = |keep[15]; // @[BFS.scala 250:125]
  wire [30:0] _select_T_48 = _select_T_46 ? 31'h8000 : 31'h0; // @[Mux.scala 98:16]
  wire [30:0] _select_T_49 = _select_T_43 ? 31'h4000 : _select_T_48; // @[Mux.scala 98:16]
  wire [30:0] _select_T_50 = _select_T_40 ? 31'h2000 : _select_T_49; // @[Mux.scala 98:16]
  wire [30:0] _select_T_51 = _select_T_37 ? 31'h1000 : _select_T_50; // @[Mux.scala 98:16]
  wire [30:0] _select_T_52 = _select_T_34 ? 31'h800 : _select_T_51; // @[Mux.scala 98:16]
  wire [30:0] _select_T_53 = _select_T_31 ? 31'h400 : _select_T_52; // @[Mux.scala 98:16]
  wire [30:0] _select_T_54 = _select_T_28 ? 31'h200 : _select_T_53; // @[Mux.scala 98:16]
  wire [30:0] _select_T_55 = _select_T_25 ? 31'h100 : _select_T_54; // @[Mux.scala 98:16]
  wire [30:0] _select_T_56 = _select_T_22 ? 31'h80 : _select_T_55; // @[Mux.scala 98:16]
  wire [30:0] _select_T_57 = _select_T_19 ? 31'h40 : _select_T_56; // @[Mux.scala 98:16]
  wire [30:0] _select_T_58 = _select_T_16 ? 31'h20 : _select_T_57; // @[Mux.scala 98:16]
  wire [30:0] _select_T_59 = _select_T_13 ? 31'h10 : _select_T_58; // @[Mux.scala 98:16]
  wire [30:0] _select_T_60 = _select_T_10 ? 31'h8 : _select_T_59; // @[Mux.scala 98:16]
  wire [30:0] _select_T_61 = _select_T_7 ? 31'h4 : _select_T_60; // @[Mux.scala 98:16]
  wire [30:0] _select_T_62 = _select_T_4 ? 31'h2 : _select_T_61; // @[Mux.scala 98:16]
  wire [30:0] select = _select_T_1 ? 31'h1 : _select_T_62; // @[Mux.scala 98:16]
  wire [31:0] _io_ddr_out_bits_tdata_T_32 = select[0] ? data[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_33 = select[1] ? data[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_34 = select[2] ? data[95:64] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_35 = select[3] ? data[127:96] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_36 = select[4] ? data[159:128] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_37 = select[5] ? data[191:160] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_38 = select[6] ? data[223:192] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_39 = select[7] ? data[255:224] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_40 = select[8] ? data[287:256] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_41 = select[9] ? data[319:288] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_42 = select[10] ? data[351:320] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_43 = select[11] ? data[383:352] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_44 = select[12] ? data[415:384] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_45 = select[13] ? data[447:416] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_46 = select[14] ? data[479:448] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_47 = select[15] ? data[511:480] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_48 = _io_ddr_out_bits_tdata_T_32 | _io_ddr_out_bits_tdata_T_33; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_49 = _io_ddr_out_bits_tdata_T_48 | _io_ddr_out_bits_tdata_T_34; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_50 = _io_ddr_out_bits_tdata_T_49 | _io_ddr_out_bits_tdata_T_35; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_51 = _io_ddr_out_bits_tdata_T_50 | _io_ddr_out_bits_tdata_T_36; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_52 = _io_ddr_out_bits_tdata_T_51 | _io_ddr_out_bits_tdata_T_37; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_53 = _io_ddr_out_bits_tdata_T_52 | _io_ddr_out_bits_tdata_T_38; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_54 = _io_ddr_out_bits_tdata_T_53 | _io_ddr_out_bits_tdata_T_39; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_55 = _io_ddr_out_bits_tdata_T_54 | _io_ddr_out_bits_tdata_T_40; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_56 = _io_ddr_out_bits_tdata_T_55 | _io_ddr_out_bits_tdata_T_41; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_57 = _io_ddr_out_bits_tdata_T_56 | _io_ddr_out_bits_tdata_T_42; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_58 = _io_ddr_out_bits_tdata_T_57 | _io_ddr_out_bits_tdata_T_43; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_59 = _io_ddr_out_bits_tdata_T_58 | _io_ddr_out_bits_tdata_T_44; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_60 = _io_ddr_out_bits_tdata_T_59 | _io_ddr_out_bits_tdata_T_45; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_61 = _io_ddr_out_bits_tdata_T_60 | _io_ddr_out_bits_tdata_T_46; // @[Mux.scala 27:72]
  wire  next_keep_0 = select[0] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_1 = select[1] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_2 = select[2] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_3 = select[3] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_4 = select[4] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_5 = select[5] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_6 = select[6] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_7 = select[7] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_8 = select[8] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_9 = select[9] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_10 = select[10] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_11 = select[11] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_12 = select[12] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_13 = select[13] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_14 = select[14] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_15 = select[15] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire [7:0] keep_lo = {next_keep_7,next_keep_6,next_keep_5,next_keep_4,next_keep_3,next_keep_2,next_keep_1,next_keep_0}
    ; // @[BFS.scala 266:36]
  wire [15:0] _keep_T = {next_keep_15,next_keep_14,next_keep_13,next_keep_12,next_keep_11,next_keep_10,next_keep_9,
    next_keep_8,keep_lo}; // @[BFS.scala 266:36]
  wire [15:0] _keep_T_1 = keep & _keep_T; // @[BFS.scala 266:18]
  assign io_xbar_in_ready = ~(|keep); // @[BFS.scala 247:23]
  assign io_ddr_out_valid = |select; // @[BFS.scala 251:33]
  assign io_ddr_out_bits_tdata = _io_ddr_out_bits_tdata_T_61 | _io_ddr_out_bits_tdata_T_47; // @[Mux.scala 27:72]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 241:21]
      data <= 512'h0; // @[BFS.scala 241:21]
    end else if (io_xbar_in_valid & io_xbar_in_ready) begin // @[BFS.scala 244:45]
      data <= io_xbar_in_bits_tdata; // @[BFS.scala 245:10]
    end
    if (reset) begin // @[BFS.scala 242:21]
      keep <= 16'h0; // @[BFS.scala 242:21]
    end else if (_T) begin // @[BFS.scala 263:45]
      keep <= io_xbar_in_bits_tkeep; // @[BFS.scala 264:10]
    end else if (io_ddr_out_valid & io_ddr_out_ready) begin // @[BFS.scala 265:52]
      keep <= _keep_T_1; // @[BFS.scala 266:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  data = _RAND_0[511:0];
  _RAND_1 = {1{`RANDOM}};
  keep = _RAND_1[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_arbitrator_17(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [127:0] io_xbar_in_bits_tdata,
  input  [3:0]   io_xbar_in_bits_tkeep,
  input          io_ddr_out_ready,
  output         io_ddr_out_valid,
  output [31:0]  io_ddr_out_bits_tdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] data; // @[BFS.scala 241:21]
  reg [3:0] keep; // @[BFS.scala 242:21]
  wire  _T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 244:25]
  wire  _select_T_1 = |keep[0]; // @[BFS.scala 250:125]
  wire  _select_T_4 = |keep[1]; // @[BFS.scala 250:125]
  wire  _select_T_7 = |keep[2]; // @[BFS.scala 250:125]
  wire  _select_T_10 = |keep[3]; // @[BFS.scala 250:125]
  wire [6:0] _select_T_12 = _select_T_10 ? 7'h8 : 7'h0; // @[Mux.scala 98:16]
  wire [6:0] _select_T_13 = _select_T_7 ? 7'h4 : _select_T_12; // @[Mux.scala 98:16]
  wire [6:0] _select_T_14 = _select_T_4 ? 7'h2 : _select_T_13; // @[Mux.scala 98:16]
  wire [6:0] select = _select_T_1 ? 7'h1 : _select_T_14; // @[Mux.scala 98:16]
  wire [31:0] _io_ddr_out_bits_tdata_T_8 = select[0] ? data[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_9 = select[1] ? data[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_10 = select[2] ? data[95:64] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_11 = select[3] ? data[127:96] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_12 = _io_ddr_out_bits_tdata_T_8 | _io_ddr_out_bits_tdata_T_9; // @[Mux.scala 27:72]
  wire [31:0] _io_ddr_out_bits_tdata_T_13 = _io_ddr_out_bits_tdata_T_12 | _io_ddr_out_bits_tdata_T_10; // @[Mux.scala 27:72]
  wire  next_keep_0 = select[0] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_1 = select[1] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_2 = select[2] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire  next_keep_3 = select[3] ? 1'h0 : 1'h1; // @[BFS.scala 261:28]
  wire [3:0] _keep_T = {next_keep_3,next_keep_2,next_keep_1,next_keep_0}; // @[BFS.scala 266:36]
  wire [3:0] _keep_T_1 = keep & _keep_T; // @[BFS.scala 266:18]
  assign io_xbar_in_ready = ~(|keep); // @[BFS.scala 247:23]
  assign io_ddr_out_valid = |select; // @[BFS.scala 251:33]
  assign io_ddr_out_bits_tdata = _io_ddr_out_bits_tdata_T_13 | _io_ddr_out_bits_tdata_T_11; // @[Mux.scala 27:72]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 241:21]
      data <= 128'h0; // @[BFS.scala 241:21]
    end else if (io_xbar_in_valid & io_xbar_in_ready) begin // @[BFS.scala 244:45]
      data <= io_xbar_in_bits_tdata; // @[BFS.scala 245:10]
    end
    if (reset) begin // @[BFS.scala 242:21]
      keep <= 4'h0; // @[BFS.scala 242:21]
    end else if (_T) begin // @[BFS.scala 263:45]
      keep <= io_xbar_in_bits_tkeep; // @[BFS.scala 264:10]
    end else if (io_ddr_out_valid & io_ddr_out_ready) begin // @[BFS.scala 265:52]
      keep <= _keep_T_1; // @[BFS.scala 266:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  data = _RAND_0[127:0];
  _RAND_1 = {1{`RANDOM}};
  keep = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Gather(
  input          clock,
  input          reset,
  output         io_ddr_in_ready,
  input          io_ddr_in_valid,
  input  [511:0] io_ddr_in_bits_tdata,
  input  [15:0]  io_ddr_in_bits_tkeep,
  input          io_gather_out_0_ready,
  output         io_gather_out_0_valid,
  output [31:0]  io_gather_out_0_bits_tdata,
  input          io_gather_out_1_ready,
  output         io_gather_out_1_valid,
  output [31:0]  io_gather_out_1_bits_tdata,
  input          io_gather_out_2_ready,
  output         io_gather_out_2_valid,
  output [31:0]  io_gather_out_2_bits_tdata,
  input          io_gather_out_3_ready,
  output         io_gather_out_3_valid,
  output [31:0]  io_gather_out_3_bits_tdata,
  input          io_gather_out_4_ready,
  output         io_gather_out_4_valid,
  output [31:0]  io_gather_out_4_bits_tdata
);
  wire  broadcaster_aclk; // @[BFS.scala 278:27]
  wire  broadcaster_aresetn; // @[BFS.scala 278:27]
  wire [511:0] broadcaster_s_axis_tdata; // @[BFS.scala 278:27]
  wire [63:0] broadcaster_s_axis_tkeep; // @[BFS.scala 278:27]
  wire  broadcaster_s_axis_tlast; // @[BFS.scala 278:27]
  wire  broadcaster_s_axis_tvalid; // @[BFS.scala 278:27]
  wire  broadcaster_s_axis_tready; // @[BFS.scala 278:27]
  wire  broadcaster_s_axis_tid; // @[BFS.scala 278:27]
  wire [2559:0] broadcaster_m_axis_tdata; // @[BFS.scala 278:27]
  wire [319:0] broadcaster_m_axis_tkeep; // @[BFS.scala 278:27]
  wire [4:0] broadcaster_m_axis_tlast; // @[BFS.scala 278:27]
  wire [4:0] broadcaster_m_axis_tvalid; // @[BFS.scala 278:27]
  wire [4:0] broadcaster_m_axis_tready; // @[BFS.scala 278:27]
  wire [4:0] broadcaster_m_axis_tid; // @[BFS.scala 278:27]
  wire  v2Apply_fifo_s_axis_aclk; // @[BFS.scala 285:28]
  wire  v2Apply_fifo_s_axis_aresetn; // @[BFS.scala 285:28]
  wire [511:0] v2Apply_fifo_s_axis_tdata; // @[BFS.scala 285:28]
  wire [63:0] v2Apply_fifo_s_axis_tkeep; // @[BFS.scala 285:28]
  wire  v2Apply_fifo_s_axis_tlast; // @[BFS.scala 285:28]
  wire  v2Apply_fifo_s_axis_tvalid; // @[BFS.scala 285:28]
  wire  v2Apply_fifo_s_axis_tready; // @[BFS.scala 285:28]
  wire  v2Apply_fifo_s_axis_tid; // @[BFS.scala 285:28]
  wire [511:0] v2Apply_fifo_m_axis_tdata; // @[BFS.scala 285:28]
  wire [63:0] v2Apply_fifo_m_axis_tkeep; // @[BFS.scala 285:28]
  wire  v2Apply_fifo_m_axis_tlast; // @[BFS.scala 285:28]
  wire  v2Apply_fifo_m_axis_tvalid; // @[BFS.scala 285:28]
  wire  v2Apply_fifo_m_axis_tready; // @[BFS.scala 285:28]
  wire  v2Apply_fifo_m_axis_tid; // @[BFS.scala 285:28]
  wire  v2Broadcast_fifo_0_s_axis_aclk; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_0_s_axis_aresetn; // @[BFS.scala 294:16]
  wire [127:0] v2Broadcast_fifo_0_s_axis_tdata; // @[BFS.scala 294:16]
  wire [15:0] v2Broadcast_fifo_0_s_axis_tkeep; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_0_s_axis_tlast; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_0_s_axis_tvalid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_0_s_axis_tready; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_0_s_axis_tid; // @[BFS.scala 294:16]
  wire [127:0] v2Broadcast_fifo_0_m_axis_tdata; // @[BFS.scala 294:16]
  wire [15:0] v2Broadcast_fifo_0_m_axis_tkeep; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_0_m_axis_tlast; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_0_m_axis_tvalid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_0_m_axis_tready; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_0_m_axis_tid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_s_axis_aclk; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_s_axis_aresetn; // @[BFS.scala 294:16]
  wire [127:0] v2Broadcast_fifo_1_s_axis_tdata; // @[BFS.scala 294:16]
  wire [15:0] v2Broadcast_fifo_1_s_axis_tkeep; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_s_axis_tlast; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_s_axis_tvalid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_s_axis_tready; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_s_axis_tid; // @[BFS.scala 294:16]
  wire [127:0] v2Broadcast_fifo_1_m_axis_tdata; // @[BFS.scala 294:16]
  wire [15:0] v2Broadcast_fifo_1_m_axis_tkeep; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_m_axis_tlast; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_m_axis_tvalid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_m_axis_tready; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_1_m_axis_tid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_s_axis_aclk; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_s_axis_aresetn; // @[BFS.scala 294:16]
  wire [127:0] v2Broadcast_fifo_2_s_axis_tdata; // @[BFS.scala 294:16]
  wire [15:0] v2Broadcast_fifo_2_s_axis_tkeep; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_s_axis_tlast; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_s_axis_tvalid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_s_axis_tready; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_s_axis_tid; // @[BFS.scala 294:16]
  wire [127:0] v2Broadcast_fifo_2_m_axis_tdata; // @[BFS.scala 294:16]
  wire [15:0] v2Broadcast_fifo_2_m_axis_tkeep; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_m_axis_tlast; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_m_axis_tvalid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_m_axis_tready; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_2_m_axis_tid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_s_axis_aclk; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_s_axis_aresetn; // @[BFS.scala 294:16]
  wire [127:0] v2Broadcast_fifo_3_s_axis_tdata; // @[BFS.scala 294:16]
  wire [15:0] v2Broadcast_fifo_3_s_axis_tkeep; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_s_axis_tlast; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_s_axis_tvalid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_s_axis_tready; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_s_axis_tid; // @[BFS.scala 294:16]
  wire [127:0] v2Broadcast_fifo_3_m_axis_tdata; // @[BFS.scala 294:16]
  wire [15:0] v2Broadcast_fifo_3_m_axis_tkeep; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_m_axis_tlast; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_m_axis_tvalid; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_m_axis_tready; // @[BFS.scala 294:16]
  wire  v2Broadcast_fifo_3_m_axis_tid; // @[BFS.scala 294:16]
  wire  v2Apply_selecter_clock; // @[BFS.scala 323:32]
  wire  v2Apply_selecter_reset; // @[BFS.scala 323:32]
  wire  v2Apply_selecter_io_xbar_in_ready; // @[BFS.scala 323:32]
  wire  v2Apply_selecter_io_xbar_in_valid; // @[BFS.scala 323:32]
  wire [511:0] v2Apply_selecter_io_xbar_in_bits_tdata; // @[BFS.scala 323:32]
  wire [15:0] v2Apply_selecter_io_xbar_in_bits_tkeep; // @[BFS.scala 323:32]
  wire  v2Apply_selecter_io_ddr_out_ready; // @[BFS.scala 323:32]
  wire  v2Apply_selecter_io_ddr_out_valid; // @[BFS.scala 323:32]
  wire [31:0] v2Apply_selecter_io_ddr_out_bits_tdata; // @[BFS.scala 323:32]
  wire  v2Broadcast_selecter_0_clock; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_0_reset; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_ready; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_0_io_xbar_in_valid; // @[BFS.scala 330:16]
  wire [127:0] v2Broadcast_selecter_0_io_xbar_in_bits_tdata; // @[BFS.scala 330:16]
  wire [3:0] v2Broadcast_selecter_0_io_xbar_in_bits_tkeep; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_0_io_ddr_out_ready; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_0_io_ddr_out_valid; // @[BFS.scala 330:16]
  wire [31:0] v2Broadcast_selecter_0_io_ddr_out_bits_tdata; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_1_clock; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_1_reset; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_ready; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_1_io_xbar_in_valid; // @[BFS.scala 330:16]
  wire [127:0] v2Broadcast_selecter_1_io_xbar_in_bits_tdata; // @[BFS.scala 330:16]
  wire [3:0] v2Broadcast_selecter_1_io_xbar_in_bits_tkeep; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_1_io_ddr_out_ready; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_1_io_ddr_out_valid; // @[BFS.scala 330:16]
  wire [31:0] v2Broadcast_selecter_1_io_ddr_out_bits_tdata; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_2_clock; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_2_reset; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_ready; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_2_io_xbar_in_valid; // @[BFS.scala 330:16]
  wire [127:0] v2Broadcast_selecter_2_io_xbar_in_bits_tdata; // @[BFS.scala 330:16]
  wire [3:0] v2Broadcast_selecter_2_io_xbar_in_bits_tkeep; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_2_io_ddr_out_ready; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_2_io_ddr_out_valid; // @[BFS.scala 330:16]
  wire [31:0] v2Broadcast_selecter_2_io_ddr_out_bits_tdata; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_3_clock; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_3_reset; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_ready; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_3_io_xbar_in_valid; // @[BFS.scala 330:16]
  wire [127:0] v2Broadcast_selecter_3_io_xbar_in_bits_tdata; // @[BFS.scala 330:16]
  wire [3:0] v2Broadcast_selecter_3_io_xbar_in_bits_tkeep; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_3_io_ddr_out_ready; // @[BFS.scala 330:16]
  wire  v2Broadcast_selecter_3_io_ddr_out_valid; // @[BFS.scala 330:16]
  wire [31:0] v2Broadcast_selecter_3_io_ddr_out_bits_tdata; // @[BFS.scala 330:16]
  wire [63:0] v2Broadcast_fifo_0_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[159:128],broadcaster_m_axis_tdata[31:0]}
    ; // @[BFS.scala 303:16]
  wire [63:0] v2Broadcast_fifo_0_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[415:384],broadcaster_m_axis_tdata[287:
    256]}; // @[BFS.scala 303:16]
  wire  _v2Broadcast_fifo_0_io_s_axis_tvalid_T_29 = broadcaster_m_axis_tkeep[0] | broadcaster_m_axis_tkeep[4] |
    broadcaster_m_axis_tkeep[8] | broadcaster_m_axis_tkeep[12]; // @[BFS.scala 313:17]
  wire [3:0] _v2Broadcast_fifo_0_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[12],broadcaster_m_axis_tkeep[8],
    broadcaster_m_axis_tkeep[4],broadcaster_m_axis_tkeep[0]}; // @[BFS.scala 316:16]
  wire [63:0] v2Broadcast_fifo_1_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[703:672],broadcaster_m_axis_tdata[575:
    544]}; // @[BFS.scala 303:16]
  wire [63:0] v2Broadcast_fifo_1_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[959:928],broadcaster_m_axis_tdata[831:
    800]}; // @[BFS.scala 303:16]
  wire  _v2Broadcast_fifo_1_io_s_axis_tvalid_T_30 = broadcaster_m_axis_tkeep[1] | broadcaster_m_axis_tkeep[5] |
    broadcaster_m_axis_tkeep[9] | broadcaster_m_axis_tkeep[13]; // @[BFS.scala 313:17]
  wire [3:0] _v2Broadcast_fifo_1_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[13],broadcaster_m_axis_tkeep[9],
    broadcaster_m_axis_tkeep[5],broadcaster_m_axis_tkeep[1]}; // @[BFS.scala 316:16]
  wire [63:0] v2Broadcast_fifo_2_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[1247:1216],broadcaster_m_axis_tdata[1119
    :1088]}; // @[BFS.scala 303:16]
  wire [63:0] v2Broadcast_fifo_2_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[1503:1472],broadcaster_m_axis_tdata[1375
    :1344]}; // @[BFS.scala 303:16]
  wire  _v2Broadcast_fifo_2_io_s_axis_tvalid_T_31 = broadcaster_m_axis_tkeep[2] | broadcaster_m_axis_tkeep[6] |
    broadcaster_m_axis_tkeep[10] | broadcaster_m_axis_tkeep[14]; // @[BFS.scala 313:17]
  wire [3:0] _v2Broadcast_fifo_2_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[14],broadcaster_m_axis_tkeep[10],
    broadcaster_m_axis_tkeep[6],broadcaster_m_axis_tkeep[2]}; // @[BFS.scala 316:16]
  wire [63:0] v2Broadcast_fifo_3_io_s_axis_tdata_lo = {broadcaster_m_axis_tdata[1791:1760],broadcaster_m_axis_tdata[1663
    :1632]}; // @[BFS.scala 303:16]
  wire [63:0] v2Broadcast_fifo_3_io_s_axis_tdata_hi = {broadcaster_m_axis_tdata[2047:2016],broadcaster_m_axis_tdata[1919
    :1888]}; // @[BFS.scala 303:16]
  wire  _v2Broadcast_fifo_3_io_s_axis_tvalid_T_32 = broadcaster_m_axis_tkeep[3] | broadcaster_m_axis_tkeep[7] |
    broadcaster_m_axis_tkeep[11] | broadcaster_m_axis_tkeep[15]; // @[BFS.scala 313:17]
  wire [3:0] _v2Broadcast_fifo_3_io_s_axis_tkeep_T_9 = {broadcaster_m_axis_tkeep[15],broadcaster_m_axis_tkeep[11],
    broadcaster_m_axis_tkeep[7],broadcaster_m_axis_tkeep[3]}; // @[BFS.scala 316:16]
  wire  _broadcaster_io_m_axis_tready_WIRE_1 = v2Broadcast_fifo_1_s_axis_tready; // @[BFS.scala 321:101 BFS.scala 321:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_0 = v2Broadcast_fifo_0_s_axis_tready; // @[BFS.scala 321:101 BFS.scala 321:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_3 = v2Broadcast_fifo_3_s_axis_tready; // @[BFS.scala 321:101 BFS.scala 321:101]
  wire  _broadcaster_io_m_axis_tready_WIRE_2 = v2Broadcast_fifo_2_s_axis_tready; // @[BFS.scala 321:101 BFS.scala 321:101]
  wire [3:0] broadcaster_io_m_axis_tready_lo_1 = {_broadcaster_io_m_axis_tready_WIRE_3,
    _broadcaster_io_m_axis_tready_WIRE_2,_broadcaster_io_m_axis_tready_WIRE_1,_broadcaster_io_m_axis_tready_WIRE_0}; // @[BFS.scala 321:151]
  wire [63:0] _v2Apply_selecter_io_xbar_in_bits_tkeep_T = v2Apply_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 124:21]
  wire [15:0] _v2Broadcast_selecter_0_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_0_m_axis_tkeep; // @[nf_arm_doce_top.scala 124:21]
  wire [15:0] _v2Broadcast_selecter_1_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_1_m_axis_tkeep; // @[nf_arm_doce_top.scala 124:21]
  wire [15:0] _v2Broadcast_selecter_2_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_2_m_axis_tkeep; // @[nf_arm_doce_top.scala 124:21]
  wire [15:0] _v2Broadcast_selecter_3_io_xbar_in_bits_tkeep_T = v2Broadcast_fifo_3_m_axis_tkeep; // @[nf_arm_doce_top.scala 124:21]
  gather_broadcaster broadcaster ( // @[BFS.scala 278:27]
    .aclk(broadcaster_aclk),
    .aresetn(broadcaster_aresetn),
    .s_axis_tdata(broadcaster_s_axis_tdata),
    .s_axis_tkeep(broadcaster_s_axis_tkeep),
    .s_axis_tlast(broadcaster_s_axis_tlast),
    .s_axis_tvalid(broadcaster_s_axis_tvalid),
    .s_axis_tready(broadcaster_s_axis_tready),
    .s_axis_tid(broadcaster_s_axis_tid),
    .m_axis_tdata(broadcaster_m_axis_tdata),
    .m_axis_tkeep(broadcaster_m_axis_tkeep),
    .m_axis_tlast(broadcaster_m_axis_tlast),
    .m_axis_tvalid(broadcaster_m_axis_tvalid),
    .m_axis_tready(broadcaster_m_axis_tready),
    .m_axis_tid(broadcaster_m_axis_tid)
  );
  v2A_fifo v2Apply_fifo ( // @[BFS.scala 285:28]
    .s_axis_aclk(v2Apply_fifo_s_axis_aclk),
    .s_axis_aresetn(v2Apply_fifo_s_axis_aresetn),
    .s_axis_tdata(v2Apply_fifo_s_axis_tdata),
    .s_axis_tkeep(v2Apply_fifo_s_axis_tkeep),
    .s_axis_tlast(v2Apply_fifo_s_axis_tlast),
    .s_axis_tvalid(v2Apply_fifo_s_axis_tvalid),
    .s_axis_tready(v2Apply_fifo_s_axis_tready),
    .s_axis_tid(v2Apply_fifo_s_axis_tid),
    .m_axis_tdata(v2Apply_fifo_m_axis_tdata),
    .m_axis_tkeep(v2Apply_fifo_m_axis_tkeep),
    .m_axis_tlast(v2Apply_fifo_m_axis_tlast),
    .m_axis_tvalid(v2Apply_fifo_m_axis_tvalid),
    .m_axis_tready(v2Apply_fifo_m_axis_tready),
    .m_axis_tid(v2Apply_fifo_m_axis_tid)
  );
  v2B_fifo v2Broadcast_fifo_0 ( // @[BFS.scala 294:16]
    .s_axis_aclk(v2Broadcast_fifo_0_s_axis_aclk),
    .s_axis_aresetn(v2Broadcast_fifo_0_s_axis_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_0_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_0_s_axis_tkeep),
    .s_axis_tlast(v2Broadcast_fifo_0_s_axis_tlast),
    .s_axis_tvalid(v2Broadcast_fifo_0_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_0_s_axis_tready),
    .s_axis_tid(v2Broadcast_fifo_0_s_axis_tid),
    .m_axis_tdata(v2Broadcast_fifo_0_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_0_m_axis_tkeep),
    .m_axis_tlast(v2Broadcast_fifo_0_m_axis_tlast),
    .m_axis_tvalid(v2Broadcast_fifo_0_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_0_m_axis_tready),
    .m_axis_tid(v2Broadcast_fifo_0_m_axis_tid)
  );
  v2B_fifo v2Broadcast_fifo_1 ( // @[BFS.scala 294:16]
    .s_axis_aclk(v2Broadcast_fifo_1_s_axis_aclk),
    .s_axis_aresetn(v2Broadcast_fifo_1_s_axis_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_1_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_1_s_axis_tkeep),
    .s_axis_tlast(v2Broadcast_fifo_1_s_axis_tlast),
    .s_axis_tvalid(v2Broadcast_fifo_1_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_1_s_axis_tready),
    .s_axis_tid(v2Broadcast_fifo_1_s_axis_tid),
    .m_axis_tdata(v2Broadcast_fifo_1_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_1_m_axis_tkeep),
    .m_axis_tlast(v2Broadcast_fifo_1_m_axis_tlast),
    .m_axis_tvalid(v2Broadcast_fifo_1_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_1_m_axis_tready),
    .m_axis_tid(v2Broadcast_fifo_1_m_axis_tid)
  );
  v2B_fifo v2Broadcast_fifo_2 ( // @[BFS.scala 294:16]
    .s_axis_aclk(v2Broadcast_fifo_2_s_axis_aclk),
    .s_axis_aresetn(v2Broadcast_fifo_2_s_axis_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_2_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_2_s_axis_tkeep),
    .s_axis_tlast(v2Broadcast_fifo_2_s_axis_tlast),
    .s_axis_tvalid(v2Broadcast_fifo_2_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_2_s_axis_tready),
    .s_axis_tid(v2Broadcast_fifo_2_s_axis_tid),
    .m_axis_tdata(v2Broadcast_fifo_2_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_2_m_axis_tkeep),
    .m_axis_tlast(v2Broadcast_fifo_2_m_axis_tlast),
    .m_axis_tvalid(v2Broadcast_fifo_2_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_2_m_axis_tready),
    .m_axis_tid(v2Broadcast_fifo_2_m_axis_tid)
  );
  v2B_fifo v2Broadcast_fifo_3 ( // @[BFS.scala 294:16]
    .s_axis_aclk(v2Broadcast_fifo_3_s_axis_aclk),
    .s_axis_aresetn(v2Broadcast_fifo_3_s_axis_aresetn),
    .s_axis_tdata(v2Broadcast_fifo_3_s_axis_tdata),
    .s_axis_tkeep(v2Broadcast_fifo_3_s_axis_tkeep),
    .s_axis_tlast(v2Broadcast_fifo_3_s_axis_tlast),
    .s_axis_tvalid(v2Broadcast_fifo_3_s_axis_tvalid),
    .s_axis_tready(v2Broadcast_fifo_3_s_axis_tready),
    .s_axis_tid(v2Broadcast_fifo_3_s_axis_tid),
    .m_axis_tdata(v2Broadcast_fifo_3_m_axis_tdata),
    .m_axis_tkeep(v2Broadcast_fifo_3_m_axis_tkeep),
    .m_axis_tlast(v2Broadcast_fifo_3_m_axis_tlast),
    .m_axis_tvalid(v2Broadcast_fifo_3_m_axis_tvalid),
    .m_axis_tready(v2Broadcast_fifo_3_m_axis_tready),
    .m_axis_tid(v2Broadcast_fifo_3_m_axis_tid)
  );
  axis_arbitrator_16 v2Apply_selecter ( // @[BFS.scala 323:32]
    .clock(v2Apply_selecter_clock),
    .reset(v2Apply_selecter_reset),
    .io_xbar_in_ready(v2Apply_selecter_io_xbar_in_ready),
    .io_xbar_in_valid(v2Apply_selecter_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Apply_selecter_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Apply_selecter_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Apply_selecter_io_ddr_out_ready),
    .io_ddr_out_valid(v2Apply_selecter_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Apply_selecter_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_17 v2Broadcast_selecter_0 ( // @[BFS.scala 330:16]
    .clock(v2Broadcast_selecter_0_clock),
    .reset(v2Broadcast_selecter_0_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_0_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_0_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Broadcast_selecter_0_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_0_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_0_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_17 v2Broadcast_selecter_1 ( // @[BFS.scala 330:16]
    .clock(v2Broadcast_selecter_1_clock),
    .reset(v2Broadcast_selecter_1_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_1_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_1_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Broadcast_selecter_1_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_1_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_1_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_17 v2Broadcast_selecter_2 ( // @[BFS.scala 330:16]
    .clock(v2Broadcast_selecter_2_clock),
    .reset(v2Broadcast_selecter_2_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_2_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_2_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Broadcast_selecter_2_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_2_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_2_io_ddr_out_bits_tdata)
  );
  axis_arbitrator_17 v2Broadcast_selecter_3 ( // @[BFS.scala 330:16]
    .clock(v2Broadcast_selecter_3_clock),
    .reset(v2Broadcast_selecter_3_reset),
    .io_xbar_in_ready(v2Broadcast_selecter_3_io_xbar_in_ready),
    .io_xbar_in_valid(v2Broadcast_selecter_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(v2Broadcast_selecter_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(v2Broadcast_selecter_3_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(v2Broadcast_selecter_3_io_ddr_out_ready),
    .io_ddr_out_valid(v2Broadcast_selecter_3_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(v2Broadcast_selecter_3_io_ddr_out_bits_tdata)
  );
  assign io_ddr_in_ready = broadcaster_s_axis_tready; // @[BFS.scala 281:19]
  assign io_gather_out_0_valid = v2Broadcast_selecter_0_io_ddr_out_valid; // @[BFS.scala 337:20]
  assign io_gather_out_0_bits_tdata = v2Broadcast_selecter_0_io_ddr_out_bits_tdata; // @[BFS.scala 337:20]
  assign io_gather_out_1_valid = v2Broadcast_selecter_1_io_ddr_out_valid; // @[BFS.scala 337:20]
  assign io_gather_out_1_bits_tdata = v2Broadcast_selecter_1_io_ddr_out_bits_tdata; // @[BFS.scala 337:20]
  assign io_gather_out_2_valid = v2Broadcast_selecter_2_io_ddr_out_valid; // @[BFS.scala 337:20]
  assign io_gather_out_2_bits_tdata = v2Broadcast_selecter_2_io_ddr_out_bits_tdata; // @[BFS.scala 337:20]
  assign io_gather_out_3_valid = v2Broadcast_selecter_3_io_ddr_out_valid; // @[BFS.scala 337:20]
  assign io_gather_out_3_bits_tdata = v2Broadcast_selecter_3_io_ddr_out_bits_tdata; // @[BFS.scala 337:20]
  assign io_gather_out_4_valid = v2Apply_selecter_io_ddr_out_valid; // @[BFS.scala 327:31]
  assign io_gather_out_4_bits_tdata = v2Apply_selecter_io_ddr_out_bits_tdata; // @[BFS.scala 327:31]
  assign broadcaster_aclk = clock; // @[BFS.scala 283:38]
  assign broadcaster_aresetn = ~reset; // @[BFS.scala 282:29]
  assign broadcaster_s_axis_tdata = io_ddr_in_bits_tdata; // @[nf_arm_doce_top.scala 116:11]
  assign broadcaster_s_axis_tkeep = {{48'd0}, io_ddr_in_bits_tkeep}; // @[nf_arm_doce_top.scala 118:11]
  assign broadcaster_s_axis_tlast = 1'h1; // @[nf_arm_doce_top.scala 117:11]
  assign broadcaster_s_axis_tvalid = io_ddr_in_valid; // @[BFS.scala 280:32]
  assign broadcaster_s_axis_tid = 1'h0;
  assign broadcaster_m_axis_tready = {v2Apply_fifo_s_axis_tready,broadcaster_io_m_axis_tready_lo_1}; // @[Cat.scala 30:58]
  assign v2Apply_fifo_s_axis_aclk = clock; // @[BFS.scala 286:46]
  assign v2Apply_fifo_s_axis_aresetn = ~reset; // @[BFS.scala 287:37]
  assign v2Apply_fifo_s_axis_tdata = broadcaster_m_axis_tdata[2559:2048]; // @[BFS.scala 288:62]
  assign v2Apply_fifo_s_axis_tkeep = broadcaster_m_axis_tkeep[319:256]; // @[BFS.scala 290:62]
  assign v2Apply_fifo_s_axis_tlast = broadcaster_m_axis_tlast[4]; // @[BFS.scala 291:62]
  assign v2Apply_fifo_s_axis_tvalid = broadcaster_m_axis_tvalid[4]; // @[BFS.scala 289:64]
  assign v2Apply_fifo_s_axis_tid = 1'h0;
  assign v2Apply_fifo_m_axis_tready = v2Apply_selecter_io_xbar_in_ready; // @[BFS.scala 325:33]
  assign v2Broadcast_fifo_0_s_axis_aclk = clock; // @[BFS.scala 299:39]
  assign v2Broadcast_fifo_0_s_axis_aresetn = ~reset; // @[BFS.scala 298:30]
  assign v2Broadcast_fifo_0_s_axis_tdata = {v2Broadcast_fifo_0_io_s_axis_tdata_hi,v2Broadcast_fifo_0_io_s_axis_tdata_lo}
    ; // @[BFS.scala 303:16]
  assign v2Broadcast_fifo_0_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_0_io_s_axis_tkeep_T_9}; // @[BFS.scala 316:16]
  assign v2Broadcast_fifo_0_s_axis_tlast = broadcaster_m_axis_tlast[0]; // @[BFS.scala 317:55]
  assign v2Broadcast_fifo_0_s_axis_tvalid = broadcaster_m_axis_tvalid[0] & _v2Broadcast_fifo_0_io_s_axis_tvalid_T_29; // @[BFS.scala 304:61]
  assign v2Broadcast_fifo_0_s_axis_tid = 1'h0;
  assign v2Broadcast_fifo_0_m_axis_tready = v2Broadcast_selecter_0_io_xbar_in_ready; // @[BFS.scala 336:44]
  assign v2Broadcast_fifo_1_s_axis_aclk = clock; // @[BFS.scala 299:39]
  assign v2Broadcast_fifo_1_s_axis_aresetn = ~reset; // @[BFS.scala 298:30]
  assign v2Broadcast_fifo_1_s_axis_tdata = {v2Broadcast_fifo_1_io_s_axis_tdata_hi,v2Broadcast_fifo_1_io_s_axis_tdata_lo}
    ; // @[BFS.scala 303:16]
  assign v2Broadcast_fifo_1_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_1_io_s_axis_tkeep_T_9}; // @[BFS.scala 316:16]
  assign v2Broadcast_fifo_1_s_axis_tlast = broadcaster_m_axis_tlast[1]; // @[BFS.scala 317:55]
  assign v2Broadcast_fifo_1_s_axis_tvalid = broadcaster_m_axis_tvalid[1] & _v2Broadcast_fifo_1_io_s_axis_tvalid_T_30; // @[BFS.scala 304:61]
  assign v2Broadcast_fifo_1_s_axis_tid = 1'h0;
  assign v2Broadcast_fifo_1_m_axis_tready = v2Broadcast_selecter_1_io_xbar_in_ready; // @[BFS.scala 336:44]
  assign v2Broadcast_fifo_2_s_axis_aclk = clock; // @[BFS.scala 299:39]
  assign v2Broadcast_fifo_2_s_axis_aresetn = ~reset; // @[BFS.scala 298:30]
  assign v2Broadcast_fifo_2_s_axis_tdata = {v2Broadcast_fifo_2_io_s_axis_tdata_hi,v2Broadcast_fifo_2_io_s_axis_tdata_lo}
    ; // @[BFS.scala 303:16]
  assign v2Broadcast_fifo_2_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_2_io_s_axis_tkeep_T_9}; // @[BFS.scala 316:16]
  assign v2Broadcast_fifo_2_s_axis_tlast = broadcaster_m_axis_tlast[2]; // @[BFS.scala 317:55]
  assign v2Broadcast_fifo_2_s_axis_tvalid = broadcaster_m_axis_tvalid[2] & _v2Broadcast_fifo_2_io_s_axis_tvalid_T_31; // @[BFS.scala 304:61]
  assign v2Broadcast_fifo_2_s_axis_tid = 1'h0;
  assign v2Broadcast_fifo_2_m_axis_tready = v2Broadcast_selecter_2_io_xbar_in_ready; // @[BFS.scala 336:44]
  assign v2Broadcast_fifo_3_s_axis_aclk = clock; // @[BFS.scala 299:39]
  assign v2Broadcast_fifo_3_s_axis_aresetn = ~reset; // @[BFS.scala 298:30]
  assign v2Broadcast_fifo_3_s_axis_tdata = {v2Broadcast_fifo_3_io_s_axis_tdata_hi,v2Broadcast_fifo_3_io_s_axis_tdata_lo}
    ; // @[BFS.scala 303:16]
  assign v2Broadcast_fifo_3_s_axis_tkeep = {{12'd0}, _v2Broadcast_fifo_3_io_s_axis_tkeep_T_9}; // @[BFS.scala 316:16]
  assign v2Broadcast_fifo_3_s_axis_tlast = broadcaster_m_axis_tlast[3]; // @[BFS.scala 317:55]
  assign v2Broadcast_fifo_3_s_axis_tvalid = broadcaster_m_axis_tvalid[3] & _v2Broadcast_fifo_3_io_s_axis_tvalid_T_32; // @[BFS.scala 304:61]
  assign v2Broadcast_fifo_3_s_axis_tid = 1'h0;
  assign v2Broadcast_fifo_3_m_axis_tready = v2Broadcast_selecter_3_io_xbar_in_ready; // @[BFS.scala 336:44]
  assign v2Apply_selecter_clock = clock;
  assign v2Apply_selecter_reset = reset;
  assign v2Apply_selecter_io_xbar_in_valid = v2Apply_fifo_m_axis_tvalid; // @[BFS.scala 324:37]
  assign v2Apply_selecter_io_xbar_in_bits_tdata = v2Apply_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 122:21]
  assign v2Apply_selecter_io_xbar_in_bits_tkeep = _v2Apply_selecter_io_xbar_in_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 124:13]
  assign v2Apply_selecter_io_ddr_out_ready = io_gather_out_4_ready; // @[BFS.scala 327:31]
  assign v2Broadcast_selecter_0_clock = clock;
  assign v2Broadcast_selecter_0_reset = reset;
  assign v2Broadcast_selecter_0_io_xbar_in_valid = v2Broadcast_fifo_0_m_axis_tvalid; // @[BFS.scala 334:26]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tdata = v2Broadcast_fifo_0_m_axis_tdata; // @[nf_arm_doce_top.scala 122:21]
  assign v2Broadcast_selecter_0_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_0_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 124:13]
  assign v2Broadcast_selecter_0_io_ddr_out_ready = io_gather_out_0_ready; // @[BFS.scala 337:20]
  assign v2Broadcast_selecter_1_clock = clock;
  assign v2Broadcast_selecter_1_reset = reset;
  assign v2Broadcast_selecter_1_io_xbar_in_valid = v2Broadcast_fifo_1_m_axis_tvalid; // @[BFS.scala 334:26]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tdata = v2Broadcast_fifo_1_m_axis_tdata; // @[nf_arm_doce_top.scala 122:21]
  assign v2Broadcast_selecter_1_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_1_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 124:13]
  assign v2Broadcast_selecter_1_io_ddr_out_ready = io_gather_out_1_ready; // @[BFS.scala 337:20]
  assign v2Broadcast_selecter_2_clock = clock;
  assign v2Broadcast_selecter_2_reset = reset;
  assign v2Broadcast_selecter_2_io_xbar_in_valid = v2Broadcast_fifo_2_m_axis_tvalid; // @[BFS.scala 334:26]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tdata = v2Broadcast_fifo_2_m_axis_tdata; // @[nf_arm_doce_top.scala 122:21]
  assign v2Broadcast_selecter_2_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_2_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 124:13]
  assign v2Broadcast_selecter_2_io_ddr_out_ready = io_gather_out_2_ready; // @[BFS.scala 337:20]
  assign v2Broadcast_selecter_3_clock = clock;
  assign v2Broadcast_selecter_3_reset = reset;
  assign v2Broadcast_selecter_3_io_xbar_in_valid = v2Broadcast_fifo_3_m_axis_tvalid; // @[BFS.scala 334:26]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tdata = v2Broadcast_fifo_3_m_axis_tdata; // @[nf_arm_doce_top.scala 122:21]
  assign v2Broadcast_selecter_3_io_xbar_in_bits_tkeep = _v2Broadcast_selecter_3_io_xbar_in_bits_tkeep_T[3:0]; // @[nf_arm_doce_top.scala 124:13]
  assign v2Broadcast_selecter_3_io_ddr_out_ready = io_gather_out_3_ready; // @[BFS.scala 337:20]
endmodule
module URAM_cluster(
  input  [17:0] io_addra,
  input         io_clka,
  input  [47:0] io_dina,
  input         io_wea,
  input  [17:0] io_addrb,
  input         io_clkb,
  output [47:0] io_doutb
);
  wire [11:0] cluster_0_addra; // @[util.scala 123:45]
  wire  cluster_0_clka; // @[util.scala 123:45]
  wire [47:0] cluster_0_dina; // @[util.scala 123:45]
  wire [47:0] cluster_0_douta; // @[util.scala 123:45]
  wire  cluster_0_ena; // @[util.scala 123:45]
  wire  cluster_0_wea; // @[util.scala 123:45]
  wire [11:0] cluster_0_addrb; // @[util.scala 123:45]
  wire  cluster_0_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_0_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_0_doutb; // @[util.scala 123:45]
  wire  cluster_0_enb; // @[util.scala 123:45]
  wire  cluster_0_web; // @[util.scala 123:45]
  wire [11:0] cluster_1_addra; // @[util.scala 123:45]
  wire  cluster_1_clka; // @[util.scala 123:45]
  wire [47:0] cluster_1_dina; // @[util.scala 123:45]
  wire [47:0] cluster_1_douta; // @[util.scala 123:45]
  wire  cluster_1_ena; // @[util.scala 123:45]
  wire  cluster_1_wea; // @[util.scala 123:45]
  wire [11:0] cluster_1_addrb; // @[util.scala 123:45]
  wire  cluster_1_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_1_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_1_doutb; // @[util.scala 123:45]
  wire  cluster_1_enb; // @[util.scala 123:45]
  wire  cluster_1_web; // @[util.scala 123:45]
  wire [11:0] cluster_2_addra; // @[util.scala 123:45]
  wire  cluster_2_clka; // @[util.scala 123:45]
  wire [47:0] cluster_2_dina; // @[util.scala 123:45]
  wire [47:0] cluster_2_douta; // @[util.scala 123:45]
  wire  cluster_2_ena; // @[util.scala 123:45]
  wire  cluster_2_wea; // @[util.scala 123:45]
  wire [11:0] cluster_2_addrb; // @[util.scala 123:45]
  wire  cluster_2_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_2_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_2_doutb; // @[util.scala 123:45]
  wire  cluster_2_enb; // @[util.scala 123:45]
  wire  cluster_2_web; // @[util.scala 123:45]
  wire [11:0] cluster_3_addra; // @[util.scala 123:45]
  wire  cluster_3_clka; // @[util.scala 123:45]
  wire [47:0] cluster_3_dina; // @[util.scala 123:45]
  wire [47:0] cluster_3_douta; // @[util.scala 123:45]
  wire  cluster_3_ena; // @[util.scala 123:45]
  wire  cluster_3_wea; // @[util.scala 123:45]
  wire [11:0] cluster_3_addrb; // @[util.scala 123:45]
  wire  cluster_3_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_3_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_3_doutb; // @[util.scala 123:45]
  wire  cluster_3_enb; // @[util.scala 123:45]
  wire  cluster_3_web; // @[util.scala 123:45]
  wire [11:0] cluster_4_addra; // @[util.scala 123:45]
  wire  cluster_4_clka; // @[util.scala 123:45]
  wire [47:0] cluster_4_dina; // @[util.scala 123:45]
  wire [47:0] cluster_4_douta; // @[util.scala 123:45]
  wire  cluster_4_ena; // @[util.scala 123:45]
  wire  cluster_4_wea; // @[util.scala 123:45]
  wire [11:0] cluster_4_addrb; // @[util.scala 123:45]
  wire  cluster_4_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_4_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_4_doutb; // @[util.scala 123:45]
  wire  cluster_4_enb; // @[util.scala 123:45]
  wire  cluster_4_web; // @[util.scala 123:45]
  wire [11:0] cluster_5_addra; // @[util.scala 123:45]
  wire  cluster_5_clka; // @[util.scala 123:45]
  wire [47:0] cluster_5_dina; // @[util.scala 123:45]
  wire [47:0] cluster_5_douta; // @[util.scala 123:45]
  wire  cluster_5_ena; // @[util.scala 123:45]
  wire  cluster_5_wea; // @[util.scala 123:45]
  wire [11:0] cluster_5_addrb; // @[util.scala 123:45]
  wire  cluster_5_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_5_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_5_doutb; // @[util.scala 123:45]
  wire  cluster_5_enb; // @[util.scala 123:45]
  wire  cluster_5_web; // @[util.scala 123:45]
  wire [11:0] cluster_6_addra; // @[util.scala 123:45]
  wire  cluster_6_clka; // @[util.scala 123:45]
  wire [47:0] cluster_6_dina; // @[util.scala 123:45]
  wire [47:0] cluster_6_douta; // @[util.scala 123:45]
  wire  cluster_6_ena; // @[util.scala 123:45]
  wire  cluster_6_wea; // @[util.scala 123:45]
  wire [11:0] cluster_6_addrb; // @[util.scala 123:45]
  wire  cluster_6_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_6_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_6_doutb; // @[util.scala 123:45]
  wire  cluster_6_enb; // @[util.scala 123:45]
  wire  cluster_6_web; // @[util.scala 123:45]
  wire [11:0] cluster_7_addra; // @[util.scala 123:45]
  wire  cluster_7_clka; // @[util.scala 123:45]
  wire [47:0] cluster_7_dina; // @[util.scala 123:45]
  wire [47:0] cluster_7_douta; // @[util.scala 123:45]
  wire  cluster_7_ena; // @[util.scala 123:45]
  wire  cluster_7_wea; // @[util.scala 123:45]
  wire [11:0] cluster_7_addrb; // @[util.scala 123:45]
  wire  cluster_7_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_7_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_7_doutb; // @[util.scala 123:45]
  wire  cluster_7_enb; // @[util.scala 123:45]
  wire  cluster_7_web; // @[util.scala 123:45]
  wire [11:0] cluster_8_addra; // @[util.scala 123:45]
  wire  cluster_8_clka; // @[util.scala 123:45]
  wire [47:0] cluster_8_dina; // @[util.scala 123:45]
  wire [47:0] cluster_8_douta; // @[util.scala 123:45]
  wire  cluster_8_ena; // @[util.scala 123:45]
  wire  cluster_8_wea; // @[util.scala 123:45]
  wire [11:0] cluster_8_addrb; // @[util.scala 123:45]
  wire  cluster_8_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_8_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_8_doutb; // @[util.scala 123:45]
  wire  cluster_8_enb; // @[util.scala 123:45]
  wire  cluster_8_web; // @[util.scala 123:45]
  wire [11:0] cluster_9_addra; // @[util.scala 123:45]
  wire  cluster_9_clka; // @[util.scala 123:45]
  wire [47:0] cluster_9_dina; // @[util.scala 123:45]
  wire [47:0] cluster_9_douta; // @[util.scala 123:45]
  wire  cluster_9_ena; // @[util.scala 123:45]
  wire  cluster_9_wea; // @[util.scala 123:45]
  wire [11:0] cluster_9_addrb; // @[util.scala 123:45]
  wire  cluster_9_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_9_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_9_doutb; // @[util.scala 123:45]
  wire  cluster_9_enb; // @[util.scala 123:45]
  wire  cluster_9_web; // @[util.scala 123:45]
  wire [11:0] cluster_10_addra; // @[util.scala 123:45]
  wire  cluster_10_clka; // @[util.scala 123:45]
  wire [47:0] cluster_10_dina; // @[util.scala 123:45]
  wire [47:0] cluster_10_douta; // @[util.scala 123:45]
  wire  cluster_10_ena; // @[util.scala 123:45]
  wire  cluster_10_wea; // @[util.scala 123:45]
  wire [11:0] cluster_10_addrb; // @[util.scala 123:45]
  wire  cluster_10_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_10_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_10_doutb; // @[util.scala 123:45]
  wire  cluster_10_enb; // @[util.scala 123:45]
  wire  cluster_10_web; // @[util.scala 123:45]
  wire [11:0] cluster_11_addra; // @[util.scala 123:45]
  wire  cluster_11_clka; // @[util.scala 123:45]
  wire [47:0] cluster_11_dina; // @[util.scala 123:45]
  wire [47:0] cluster_11_douta; // @[util.scala 123:45]
  wire  cluster_11_ena; // @[util.scala 123:45]
  wire  cluster_11_wea; // @[util.scala 123:45]
  wire [11:0] cluster_11_addrb; // @[util.scala 123:45]
  wire  cluster_11_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_11_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_11_doutb; // @[util.scala 123:45]
  wire  cluster_11_enb; // @[util.scala 123:45]
  wire  cluster_11_web; // @[util.scala 123:45]
  wire [11:0] cluster_12_addra; // @[util.scala 123:45]
  wire  cluster_12_clka; // @[util.scala 123:45]
  wire [47:0] cluster_12_dina; // @[util.scala 123:45]
  wire [47:0] cluster_12_douta; // @[util.scala 123:45]
  wire  cluster_12_ena; // @[util.scala 123:45]
  wire  cluster_12_wea; // @[util.scala 123:45]
  wire [11:0] cluster_12_addrb; // @[util.scala 123:45]
  wire  cluster_12_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_12_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_12_doutb; // @[util.scala 123:45]
  wire  cluster_12_enb; // @[util.scala 123:45]
  wire  cluster_12_web; // @[util.scala 123:45]
  wire [11:0] cluster_13_addra; // @[util.scala 123:45]
  wire  cluster_13_clka; // @[util.scala 123:45]
  wire [47:0] cluster_13_dina; // @[util.scala 123:45]
  wire [47:0] cluster_13_douta; // @[util.scala 123:45]
  wire  cluster_13_ena; // @[util.scala 123:45]
  wire  cluster_13_wea; // @[util.scala 123:45]
  wire [11:0] cluster_13_addrb; // @[util.scala 123:45]
  wire  cluster_13_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_13_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_13_doutb; // @[util.scala 123:45]
  wire  cluster_13_enb; // @[util.scala 123:45]
  wire  cluster_13_web; // @[util.scala 123:45]
  wire [11:0] cluster_14_addra; // @[util.scala 123:45]
  wire  cluster_14_clka; // @[util.scala 123:45]
  wire [47:0] cluster_14_dina; // @[util.scala 123:45]
  wire [47:0] cluster_14_douta; // @[util.scala 123:45]
  wire  cluster_14_ena; // @[util.scala 123:45]
  wire  cluster_14_wea; // @[util.scala 123:45]
  wire [11:0] cluster_14_addrb; // @[util.scala 123:45]
  wire  cluster_14_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_14_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_14_doutb; // @[util.scala 123:45]
  wire  cluster_14_enb; // @[util.scala 123:45]
  wire  cluster_14_web; // @[util.scala 123:45]
  wire [11:0] cluster_15_addra; // @[util.scala 123:45]
  wire  cluster_15_clka; // @[util.scala 123:45]
  wire [47:0] cluster_15_dina; // @[util.scala 123:45]
  wire [47:0] cluster_15_douta; // @[util.scala 123:45]
  wire  cluster_15_ena; // @[util.scala 123:45]
  wire  cluster_15_wea; // @[util.scala 123:45]
  wire [11:0] cluster_15_addrb; // @[util.scala 123:45]
  wire  cluster_15_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_15_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_15_doutb; // @[util.scala 123:45]
  wire  cluster_15_enb; // @[util.scala 123:45]
  wire  cluster_15_web; // @[util.scala 123:45]
  wire [11:0] cluster_16_addra; // @[util.scala 123:45]
  wire  cluster_16_clka; // @[util.scala 123:45]
  wire [47:0] cluster_16_dina; // @[util.scala 123:45]
  wire [47:0] cluster_16_douta; // @[util.scala 123:45]
  wire  cluster_16_ena; // @[util.scala 123:45]
  wire  cluster_16_wea; // @[util.scala 123:45]
  wire [11:0] cluster_16_addrb; // @[util.scala 123:45]
  wire  cluster_16_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_16_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_16_doutb; // @[util.scala 123:45]
  wire  cluster_16_enb; // @[util.scala 123:45]
  wire  cluster_16_web; // @[util.scala 123:45]
  wire [11:0] cluster_17_addra; // @[util.scala 123:45]
  wire  cluster_17_clka; // @[util.scala 123:45]
  wire [47:0] cluster_17_dina; // @[util.scala 123:45]
  wire [47:0] cluster_17_douta; // @[util.scala 123:45]
  wire  cluster_17_ena; // @[util.scala 123:45]
  wire  cluster_17_wea; // @[util.scala 123:45]
  wire [11:0] cluster_17_addrb; // @[util.scala 123:45]
  wire  cluster_17_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_17_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_17_doutb; // @[util.scala 123:45]
  wire  cluster_17_enb; // @[util.scala 123:45]
  wire  cluster_17_web; // @[util.scala 123:45]
  wire [11:0] cluster_18_addra; // @[util.scala 123:45]
  wire  cluster_18_clka; // @[util.scala 123:45]
  wire [47:0] cluster_18_dina; // @[util.scala 123:45]
  wire [47:0] cluster_18_douta; // @[util.scala 123:45]
  wire  cluster_18_ena; // @[util.scala 123:45]
  wire  cluster_18_wea; // @[util.scala 123:45]
  wire [11:0] cluster_18_addrb; // @[util.scala 123:45]
  wire  cluster_18_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_18_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_18_doutb; // @[util.scala 123:45]
  wire  cluster_18_enb; // @[util.scala 123:45]
  wire  cluster_18_web; // @[util.scala 123:45]
  wire [11:0] cluster_19_addra; // @[util.scala 123:45]
  wire  cluster_19_clka; // @[util.scala 123:45]
  wire [47:0] cluster_19_dina; // @[util.scala 123:45]
  wire [47:0] cluster_19_douta; // @[util.scala 123:45]
  wire  cluster_19_ena; // @[util.scala 123:45]
  wire  cluster_19_wea; // @[util.scala 123:45]
  wire [11:0] cluster_19_addrb; // @[util.scala 123:45]
  wire  cluster_19_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_19_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_19_doutb; // @[util.scala 123:45]
  wire  cluster_19_enb; // @[util.scala 123:45]
  wire  cluster_19_web; // @[util.scala 123:45]
  wire [11:0] cluster_20_addra; // @[util.scala 123:45]
  wire  cluster_20_clka; // @[util.scala 123:45]
  wire [47:0] cluster_20_dina; // @[util.scala 123:45]
  wire [47:0] cluster_20_douta; // @[util.scala 123:45]
  wire  cluster_20_ena; // @[util.scala 123:45]
  wire  cluster_20_wea; // @[util.scala 123:45]
  wire [11:0] cluster_20_addrb; // @[util.scala 123:45]
  wire  cluster_20_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_20_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_20_doutb; // @[util.scala 123:45]
  wire  cluster_20_enb; // @[util.scala 123:45]
  wire  cluster_20_web; // @[util.scala 123:45]
  wire [11:0] cluster_21_addra; // @[util.scala 123:45]
  wire  cluster_21_clka; // @[util.scala 123:45]
  wire [47:0] cluster_21_dina; // @[util.scala 123:45]
  wire [47:0] cluster_21_douta; // @[util.scala 123:45]
  wire  cluster_21_ena; // @[util.scala 123:45]
  wire  cluster_21_wea; // @[util.scala 123:45]
  wire [11:0] cluster_21_addrb; // @[util.scala 123:45]
  wire  cluster_21_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_21_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_21_doutb; // @[util.scala 123:45]
  wire  cluster_21_enb; // @[util.scala 123:45]
  wire  cluster_21_web; // @[util.scala 123:45]
  wire [11:0] cluster_22_addra; // @[util.scala 123:45]
  wire  cluster_22_clka; // @[util.scala 123:45]
  wire [47:0] cluster_22_dina; // @[util.scala 123:45]
  wire [47:0] cluster_22_douta; // @[util.scala 123:45]
  wire  cluster_22_ena; // @[util.scala 123:45]
  wire  cluster_22_wea; // @[util.scala 123:45]
  wire [11:0] cluster_22_addrb; // @[util.scala 123:45]
  wire  cluster_22_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_22_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_22_doutb; // @[util.scala 123:45]
  wire  cluster_22_enb; // @[util.scala 123:45]
  wire  cluster_22_web; // @[util.scala 123:45]
  wire [11:0] cluster_23_addra; // @[util.scala 123:45]
  wire  cluster_23_clka; // @[util.scala 123:45]
  wire [47:0] cluster_23_dina; // @[util.scala 123:45]
  wire [47:0] cluster_23_douta; // @[util.scala 123:45]
  wire  cluster_23_ena; // @[util.scala 123:45]
  wire  cluster_23_wea; // @[util.scala 123:45]
  wire [11:0] cluster_23_addrb; // @[util.scala 123:45]
  wire  cluster_23_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_23_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_23_doutb; // @[util.scala 123:45]
  wire  cluster_23_enb; // @[util.scala 123:45]
  wire  cluster_23_web; // @[util.scala 123:45]
  wire [11:0] cluster_24_addra; // @[util.scala 123:45]
  wire  cluster_24_clka; // @[util.scala 123:45]
  wire [47:0] cluster_24_dina; // @[util.scala 123:45]
  wire [47:0] cluster_24_douta; // @[util.scala 123:45]
  wire  cluster_24_ena; // @[util.scala 123:45]
  wire  cluster_24_wea; // @[util.scala 123:45]
  wire [11:0] cluster_24_addrb; // @[util.scala 123:45]
  wire  cluster_24_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_24_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_24_doutb; // @[util.scala 123:45]
  wire  cluster_24_enb; // @[util.scala 123:45]
  wire  cluster_24_web; // @[util.scala 123:45]
  wire [11:0] cluster_25_addra; // @[util.scala 123:45]
  wire  cluster_25_clka; // @[util.scala 123:45]
  wire [47:0] cluster_25_dina; // @[util.scala 123:45]
  wire [47:0] cluster_25_douta; // @[util.scala 123:45]
  wire  cluster_25_ena; // @[util.scala 123:45]
  wire  cluster_25_wea; // @[util.scala 123:45]
  wire [11:0] cluster_25_addrb; // @[util.scala 123:45]
  wire  cluster_25_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_25_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_25_doutb; // @[util.scala 123:45]
  wire  cluster_25_enb; // @[util.scala 123:45]
  wire  cluster_25_web; // @[util.scala 123:45]
  wire [11:0] cluster_26_addra; // @[util.scala 123:45]
  wire  cluster_26_clka; // @[util.scala 123:45]
  wire [47:0] cluster_26_dina; // @[util.scala 123:45]
  wire [47:0] cluster_26_douta; // @[util.scala 123:45]
  wire  cluster_26_ena; // @[util.scala 123:45]
  wire  cluster_26_wea; // @[util.scala 123:45]
  wire [11:0] cluster_26_addrb; // @[util.scala 123:45]
  wire  cluster_26_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_26_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_26_doutb; // @[util.scala 123:45]
  wire  cluster_26_enb; // @[util.scala 123:45]
  wire  cluster_26_web; // @[util.scala 123:45]
  wire [11:0] cluster_27_addra; // @[util.scala 123:45]
  wire  cluster_27_clka; // @[util.scala 123:45]
  wire [47:0] cluster_27_dina; // @[util.scala 123:45]
  wire [47:0] cluster_27_douta; // @[util.scala 123:45]
  wire  cluster_27_ena; // @[util.scala 123:45]
  wire  cluster_27_wea; // @[util.scala 123:45]
  wire [11:0] cluster_27_addrb; // @[util.scala 123:45]
  wire  cluster_27_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_27_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_27_doutb; // @[util.scala 123:45]
  wire  cluster_27_enb; // @[util.scala 123:45]
  wire  cluster_27_web; // @[util.scala 123:45]
  wire [11:0] cluster_28_addra; // @[util.scala 123:45]
  wire  cluster_28_clka; // @[util.scala 123:45]
  wire [47:0] cluster_28_dina; // @[util.scala 123:45]
  wire [47:0] cluster_28_douta; // @[util.scala 123:45]
  wire  cluster_28_ena; // @[util.scala 123:45]
  wire  cluster_28_wea; // @[util.scala 123:45]
  wire [11:0] cluster_28_addrb; // @[util.scala 123:45]
  wire  cluster_28_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_28_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_28_doutb; // @[util.scala 123:45]
  wire  cluster_28_enb; // @[util.scala 123:45]
  wire  cluster_28_web; // @[util.scala 123:45]
  wire [11:0] cluster_29_addra; // @[util.scala 123:45]
  wire  cluster_29_clka; // @[util.scala 123:45]
  wire [47:0] cluster_29_dina; // @[util.scala 123:45]
  wire [47:0] cluster_29_douta; // @[util.scala 123:45]
  wire  cluster_29_ena; // @[util.scala 123:45]
  wire  cluster_29_wea; // @[util.scala 123:45]
  wire [11:0] cluster_29_addrb; // @[util.scala 123:45]
  wire  cluster_29_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_29_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_29_doutb; // @[util.scala 123:45]
  wire  cluster_29_enb; // @[util.scala 123:45]
  wire  cluster_29_web; // @[util.scala 123:45]
  wire [11:0] cluster_30_addra; // @[util.scala 123:45]
  wire  cluster_30_clka; // @[util.scala 123:45]
  wire [47:0] cluster_30_dina; // @[util.scala 123:45]
  wire [47:0] cluster_30_douta; // @[util.scala 123:45]
  wire  cluster_30_ena; // @[util.scala 123:45]
  wire  cluster_30_wea; // @[util.scala 123:45]
  wire [11:0] cluster_30_addrb; // @[util.scala 123:45]
  wire  cluster_30_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_30_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_30_doutb; // @[util.scala 123:45]
  wire  cluster_30_enb; // @[util.scala 123:45]
  wire  cluster_30_web; // @[util.scala 123:45]
  wire [11:0] cluster_31_addra; // @[util.scala 123:45]
  wire  cluster_31_clka; // @[util.scala 123:45]
  wire [47:0] cluster_31_dina; // @[util.scala 123:45]
  wire [47:0] cluster_31_douta; // @[util.scala 123:45]
  wire  cluster_31_ena; // @[util.scala 123:45]
  wire  cluster_31_wea; // @[util.scala 123:45]
  wire [11:0] cluster_31_addrb; // @[util.scala 123:45]
  wire  cluster_31_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_31_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_31_doutb; // @[util.scala 123:45]
  wire  cluster_31_enb; // @[util.scala 123:45]
  wire  cluster_31_web; // @[util.scala 123:45]
  wire [11:0] cluster_32_addra; // @[util.scala 123:45]
  wire  cluster_32_clka; // @[util.scala 123:45]
  wire [47:0] cluster_32_dina; // @[util.scala 123:45]
  wire [47:0] cluster_32_douta; // @[util.scala 123:45]
  wire  cluster_32_ena; // @[util.scala 123:45]
  wire  cluster_32_wea; // @[util.scala 123:45]
  wire [11:0] cluster_32_addrb; // @[util.scala 123:45]
  wire  cluster_32_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_32_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_32_doutb; // @[util.scala 123:45]
  wire  cluster_32_enb; // @[util.scala 123:45]
  wire  cluster_32_web; // @[util.scala 123:45]
  wire [11:0] cluster_33_addra; // @[util.scala 123:45]
  wire  cluster_33_clka; // @[util.scala 123:45]
  wire [47:0] cluster_33_dina; // @[util.scala 123:45]
  wire [47:0] cluster_33_douta; // @[util.scala 123:45]
  wire  cluster_33_ena; // @[util.scala 123:45]
  wire  cluster_33_wea; // @[util.scala 123:45]
  wire [11:0] cluster_33_addrb; // @[util.scala 123:45]
  wire  cluster_33_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_33_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_33_doutb; // @[util.scala 123:45]
  wire  cluster_33_enb; // @[util.scala 123:45]
  wire  cluster_33_web; // @[util.scala 123:45]
  wire [11:0] cluster_34_addra; // @[util.scala 123:45]
  wire  cluster_34_clka; // @[util.scala 123:45]
  wire [47:0] cluster_34_dina; // @[util.scala 123:45]
  wire [47:0] cluster_34_douta; // @[util.scala 123:45]
  wire  cluster_34_ena; // @[util.scala 123:45]
  wire  cluster_34_wea; // @[util.scala 123:45]
  wire [11:0] cluster_34_addrb; // @[util.scala 123:45]
  wire  cluster_34_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_34_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_34_doutb; // @[util.scala 123:45]
  wire  cluster_34_enb; // @[util.scala 123:45]
  wire  cluster_34_web; // @[util.scala 123:45]
  wire [11:0] cluster_35_addra; // @[util.scala 123:45]
  wire  cluster_35_clka; // @[util.scala 123:45]
  wire [47:0] cluster_35_dina; // @[util.scala 123:45]
  wire [47:0] cluster_35_douta; // @[util.scala 123:45]
  wire  cluster_35_ena; // @[util.scala 123:45]
  wire  cluster_35_wea; // @[util.scala 123:45]
  wire [11:0] cluster_35_addrb; // @[util.scala 123:45]
  wire  cluster_35_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_35_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_35_doutb; // @[util.scala 123:45]
  wire  cluster_35_enb; // @[util.scala 123:45]
  wire  cluster_35_web; // @[util.scala 123:45]
  wire [11:0] cluster_36_addra; // @[util.scala 123:45]
  wire  cluster_36_clka; // @[util.scala 123:45]
  wire [47:0] cluster_36_dina; // @[util.scala 123:45]
  wire [47:0] cluster_36_douta; // @[util.scala 123:45]
  wire  cluster_36_ena; // @[util.scala 123:45]
  wire  cluster_36_wea; // @[util.scala 123:45]
  wire [11:0] cluster_36_addrb; // @[util.scala 123:45]
  wire  cluster_36_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_36_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_36_doutb; // @[util.scala 123:45]
  wire  cluster_36_enb; // @[util.scala 123:45]
  wire  cluster_36_web; // @[util.scala 123:45]
  wire [11:0] cluster_37_addra; // @[util.scala 123:45]
  wire  cluster_37_clka; // @[util.scala 123:45]
  wire [47:0] cluster_37_dina; // @[util.scala 123:45]
  wire [47:0] cluster_37_douta; // @[util.scala 123:45]
  wire  cluster_37_ena; // @[util.scala 123:45]
  wire  cluster_37_wea; // @[util.scala 123:45]
  wire [11:0] cluster_37_addrb; // @[util.scala 123:45]
  wire  cluster_37_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_37_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_37_doutb; // @[util.scala 123:45]
  wire  cluster_37_enb; // @[util.scala 123:45]
  wire  cluster_37_web; // @[util.scala 123:45]
  wire [11:0] cluster_38_addra; // @[util.scala 123:45]
  wire  cluster_38_clka; // @[util.scala 123:45]
  wire [47:0] cluster_38_dina; // @[util.scala 123:45]
  wire [47:0] cluster_38_douta; // @[util.scala 123:45]
  wire  cluster_38_ena; // @[util.scala 123:45]
  wire  cluster_38_wea; // @[util.scala 123:45]
  wire [11:0] cluster_38_addrb; // @[util.scala 123:45]
  wire  cluster_38_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_38_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_38_doutb; // @[util.scala 123:45]
  wire  cluster_38_enb; // @[util.scala 123:45]
  wire  cluster_38_web; // @[util.scala 123:45]
  wire [11:0] cluster_39_addra; // @[util.scala 123:45]
  wire  cluster_39_clka; // @[util.scala 123:45]
  wire [47:0] cluster_39_dina; // @[util.scala 123:45]
  wire [47:0] cluster_39_douta; // @[util.scala 123:45]
  wire  cluster_39_ena; // @[util.scala 123:45]
  wire  cluster_39_wea; // @[util.scala 123:45]
  wire [11:0] cluster_39_addrb; // @[util.scala 123:45]
  wire  cluster_39_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_39_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_39_doutb; // @[util.scala 123:45]
  wire  cluster_39_enb; // @[util.scala 123:45]
  wire  cluster_39_web; // @[util.scala 123:45]
  wire [11:0] cluster_40_addra; // @[util.scala 123:45]
  wire  cluster_40_clka; // @[util.scala 123:45]
  wire [47:0] cluster_40_dina; // @[util.scala 123:45]
  wire [47:0] cluster_40_douta; // @[util.scala 123:45]
  wire  cluster_40_ena; // @[util.scala 123:45]
  wire  cluster_40_wea; // @[util.scala 123:45]
  wire [11:0] cluster_40_addrb; // @[util.scala 123:45]
  wire  cluster_40_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_40_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_40_doutb; // @[util.scala 123:45]
  wire  cluster_40_enb; // @[util.scala 123:45]
  wire  cluster_40_web; // @[util.scala 123:45]
  wire [11:0] cluster_41_addra; // @[util.scala 123:45]
  wire  cluster_41_clka; // @[util.scala 123:45]
  wire [47:0] cluster_41_dina; // @[util.scala 123:45]
  wire [47:0] cluster_41_douta; // @[util.scala 123:45]
  wire  cluster_41_ena; // @[util.scala 123:45]
  wire  cluster_41_wea; // @[util.scala 123:45]
  wire [11:0] cluster_41_addrb; // @[util.scala 123:45]
  wire  cluster_41_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_41_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_41_doutb; // @[util.scala 123:45]
  wire  cluster_41_enb; // @[util.scala 123:45]
  wire  cluster_41_web; // @[util.scala 123:45]
  wire [11:0] cluster_42_addra; // @[util.scala 123:45]
  wire  cluster_42_clka; // @[util.scala 123:45]
  wire [47:0] cluster_42_dina; // @[util.scala 123:45]
  wire [47:0] cluster_42_douta; // @[util.scala 123:45]
  wire  cluster_42_ena; // @[util.scala 123:45]
  wire  cluster_42_wea; // @[util.scala 123:45]
  wire [11:0] cluster_42_addrb; // @[util.scala 123:45]
  wire  cluster_42_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_42_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_42_doutb; // @[util.scala 123:45]
  wire  cluster_42_enb; // @[util.scala 123:45]
  wire  cluster_42_web; // @[util.scala 123:45]
  wire [11:0] cluster_43_addra; // @[util.scala 123:45]
  wire  cluster_43_clka; // @[util.scala 123:45]
  wire [47:0] cluster_43_dina; // @[util.scala 123:45]
  wire [47:0] cluster_43_douta; // @[util.scala 123:45]
  wire  cluster_43_ena; // @[util.scala 123:45]
  wire  cluster_43_wea; // @[util.scala 123:45]
  wire [11:0] cluster_43_addrb; // @[util.scala 123:45]
  wire  cluster_43_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_43_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_43_doutb; // @[util.scala 123:45]
  wire  cluster_43_enb; // @[util.scala 123:45]
  wire  cluster_43_web; // @[util.scala 123:45]
  wire [11:0] cluster_44_addra; // @[util.scala 123:45]
  wire  cluster_44_clka; // @[util.scala 123:45]
  wire [47:0] cluster_44_dina; // @[util.scala 123:45]
  wire [47:0] cluster_44_douta; // @[util.scala 123:45]
  wire  cluster_44_ena; // @[util.scala 123:45]
  wire  cluster_44_wea; // @[util.scala 123:45]
  wire [11:0] cluster_44_addrb; // @[util.scala 123:45]
  wire  cluster_44_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_44_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_44_doutb; // @[util.scala 123:45]
  wire  cluster_44_enb; // @[util.scala 123:45]
  wire  cluster_44_web; // @[util.scala 123:45]
  wire [11:0] cluster_45_addra; // @[util.scala 123:45]
  wire  cluster_45_clka; // @[util.scala 123:45]
  wire [47:0] cluster_45_dina; // @[util.scala 123:45]
  wire [47:0] cluster_45_douta; // @[util.scala 123:45]
  wire  cluster_45_ena; // @[util.scala 123:45]
  wire  cluster_45_wea; // @[util.scala 123:45]
  wire [11:0] cluster_45_addrb; // @[util.scala 123:45]
  wire  cluster_45_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_45_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_45_doutb; // @[util.scala 123:45]
  wire  cluster_45_enb; // @[util.scala 123:45]
  wire  cluster_45_web; // @[util.scala 123:45]
  wire [11:0] cluster_46_addra; // @[util.scala 123:45]
  wire  cluster_46_clka; // @[util.scala 123:45]
  wire [47:0] cluster_46_dina; // @[util.scala 123:45]
  wire [47:0] cluster_46_douta; // @[util.scala 123:45]
  wire  cluster_46_ena; // @[util.scala 123:45]
  wire  cluster_46_wea; // @[util.scala 123:45]
  wire [11:0] cluster_46_addrb; // @[util.scala 123:45]
  wire  cluster_46_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_46_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_46_doutb; // @[util.scala 123:45]
  wire  cluster_46_enb; // @[util.scala 123:45]
  wire  cluster_46_web; // @[util.scala 123:45]
  wire [11:0] cluster_47_addra; // @[util.scala 123:45]
  wire  cluster_47_clka; // @[util.scala 123:45]
  wire [47:0] cluster_47_dina; // @[util.scala 123:45]
  wire [47:0] cluster_47_douta; // @[util.scala 123:45]
  wire  cluster_47_ena; // @[util.scala 123:45]
  wire  cluster_47_wea; // @[util.scala 123:45]
  wire [11:0] cluster_47_addrb; // @[util.scala 123:45]
  wire  cluster_47_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_47_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_47_doutb; // @[util.scala 123:45]
  wire  cluster_47_enb; // @[util.scala 123:45]
  wire  cluster_47_web; // @[util.scala 123:45]
  wire [11:0] cluster_48_addra; // @[util.scala 123:45]
  wire  cluster_48_clka; // @[util.scala 123:45]
  wire [47:0] cluster_48_dina; // @[util.scala 123:45]
  wire [47:0] cluster_48_douta; // @[util.scala 123:45]
  wire  cluster_48_ena; // @[util.scala 123:45]
  wire  cluster_48_wea; // @[util.scala 123:45]
  wire [11:0] cluster_48_addrb; // @[util.scala 123:45]
  wire  cluster_48_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_48_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_48_doutb; // @[util.scala 123:45]
  wire  cluster_48_enb; // @[util.scala 123:45]
  wire  cluster_48_web; // @[util.scala 123:45]
  wire [11:0] cluster_49_addra; // @[util.scala 123:45]
  wire  cluster_49_clka; // @[util.scala 123:45]
  wire [47:0] cluster_49_dina; // @[util.scala 123:45]
  wire [47:0] cluster_49_douta; // @[util.scala 123:45]
  wire  cluster_49_ena; // @[util.scala 123:45]
  wire  cluster_49_wea; // @[util.scala 123:45]
  wire [11:0] cluster_49_addrb; // @[util.scala 123:45]
  wire  cluster_49_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_49_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_49_doutb; // @[util.scala 123:45]
  wire  cluster_49_enb; // @[util.scala 123:45]
  wire  cluster_49_web; // @[util.scala 123:45]
  wire [11:0] cluster_50_addra; // @[util.scala 123:45]
  wire  cluster_50_clka; // @[util.scala 123:45]
  wire [47:0] cluster_50_dina; // @[util.scala 123:45]
  wire [47:0] cluster_50_douta; // @[util.scala 123:45]
  wire  cluster_50_ena; // @[util.scala 123:45]
  wire  cluster_50_wea; // @[util.scala 123:45]
  wire [11:0] cluster_50_addrb; // @[util.scala 123:45]
  wire  cluster_50_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_50_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_50_doutb; // @[util.scala 123:45]
  wire  cluster_50_enb; // @[util.scala 123:45]
  wire  cluster_50_web; // @[util.scala 123:45]
  wire [11:0] cluster_51_addra; // @[util.scala 123:45]
  wire  cluster_51_clka; // @[util.scala 123:45]
  wire [47:0] cluster_51_dina; // @[util.scala 123:45]
  wire [47:0] cluster_51_douta; // @[util.scala 123:45]
  wire  cluster_51_ena; // @[util.scala 123:45]
  wire  cluster_51_wea; // @[util.scala 123:45]
  wire [11:0] cluster_51_addrb; // @[util.scala 123:45]
  wire  cluster_51_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_51_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_51_doutb; // @[util.scala 123:45]
  wire  cluster_51_enb; // @[util.scala 123:45]
  wire  cluster_51_web; // @[util.scala 123:45]
  wire [11:0] cluster_52_addra; // @[util.scala 123:45]
  wire  cluster_52_clka; // @[util.scala 123:45]
  wire [47:0] cluster_52_dina; // @[util.scala 123:45]
  wire [47:0] cluster_52_douta; // @[util.scala 123:45]
  wire  cluster_52_ena; // @[util.scala 123:45]
  wire  cluster_52_wea; // @[util.scala 123:45]
  wire [11:0] cluster_52_addrb; // @[util.scala 123:45]
  wire  cluster_52_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_52_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_52_doutb; // @[util.scala 123:45]
  wire  cluster_52_enb; // @[util.scala 123:45]
  wire  cluster_52_web; // @[util.scala 123:45]
  wire [11:0] cluster_53_addra; // @[util.scala 123:45]
  wire  cluster_53_clka; // @[util.scala 123:45]
  wire [47:0] cluster_53_dina; // @[util.scala 123:45]
  wire [47:0] cluster_53_douta; // @[util.scala 123:45]
  wire  cluster_53_ena; // @[util.scala 123:45]
  wire  cluster_53_wea; // @[util.scala 123:45]
  wire [11:0] cluster_53_addrb; // @[util.scala 123:45]
  wire  cluster_53_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_53_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_53_doutb; // @[util.scala 123:45]
  wire  cluster_53_enb; // @[util.scala 123:45]
  wire  cluster_53_web; // @[util.scala 123:45]
  wire [11:0] cluster_54_addra; // @[util.scala 123:45]
  wire  cluster_54_clka; // @[util.scala 123:45]
  wire [47:0] cluster_54_dina; // @[util.scala 123:45]
  wire [47:0] cluster_54_douta; // @[util.scala 123:45]
  wire  cluster_54_ena; // @[util.scala 123:45]
  wire  cluster_54_wea; // @[util.scala 123:45]
  wire [11:0] cluster_54_addrb; // @[util.scala 123:45]
  wire  cluster_54_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_54_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_54_doutb; // @[util.scala 123:45]
  wire  cluster_54_enb; // @[util.scala 123:45]
  wire  cluster_54_web; // @[util.scala 123:45]
  wire [11:0] cluster_55_addra; // @[util.scala 123:45]
  wire  cluster_55_clka; // @[util.scala 123:45]
  wire [47:0] cluster_55_dina; // @[util.scala 123:45]
  wire [47:0] cluster_55_douta; // @[util.scala 123:45]
  wire  cluster_55_ena; // @[util.scala 123:45]
  wire  cluster_55_wea; // @[util.scala 123:45]
  wire [11:0] cluster_55_addrb; // @[util.scala 123:45]
  wire  cluster_55_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_55_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_55_doutb; // @[util.scala 123:45]
  wire  cluster_55_enb; // @[util.scala 123:45]
  wire  cluster_55_web; // @[util.scala 123:45]
  wire [11:0] cluster_56_addra; // @[util.scala 123:45]
  wire  cluster_56_clka; // @[util.scala 123:45]
  wire [47:0] cluster_56_dina; // @[util.scala 123:45]
  wire [47:0] cluster_56_douta; // @[util.scala 123:45]
  wire  cluster_56_ena; // @[util.scala 123:45]
  wire  cluster_56_wea; // @[util.scala 123:45]
  wire [11:0] cluster_56_addrb; // @[util.scala 123:45]
  wire  cluster_56_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_56_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_56_doutb; // @[util.scala 123:45]
  wire  cluster_56_enb; // @[util.scala 123:45]
  wire  cluster_56_web; // @[util.scala 123:45]
  wire [11:0] cluster_57_addra; // @[util.scala 123:45]
  wire  cluster_57_clka; // @[util.scala 123:45]
  wire [47:0] cluster_57_dina; // @[util.scala 123:45]
  wire [47:0] cluster_57_douta; // @[util.scala 123:45]
  wire  cluster_57_ena; // @[util.scala 123:45]
  wire  cluster_57_wea; // @[util.scala 123:45]
  wire [11:0] cluster_57_addrb; // @[util.scala 123:45]
  wire  cluster_57_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_57_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_57_doutb; // @[util.scala 123:45]
  wire  cluster_57_enb; // @[util.scala 123:45]
  wire  cluster_57_web; // @[util.scala 123:45]
  wire [11:0] cluster_58_addra; // @[util.scala 123:45]
  wire  cluster_58_clka; // @[util.scala 123:45]
  wire [47:0] cluster_58_dina; // @[util.scala 123:45]
  wire [47:0] cluster_58_douta; // @[util.scala 123:45]
  wire  cluster_58_ena; // @[util.scala 123:45]
  wire  cluster_58_wea; // @[util.scala 123:45]
  wire [11:0] cluster_58_addrb; // @[util.scala 123:45]
  wire  cluster_58_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_58_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_58_doutb; // @[util.scala 123:45]
  wire  cluster_58_enb; // @[util.scala 123:45]
  wire  cluster_58_web; // @[util.scala 123:45]
  wire [11:0] cluster_59_addra; // @[util.scala 123:45]
  wire  cluster_59_clka; // @[util.scala 123:45]
  wire [47:0] cluster_59_dina; // @[util.scala 123:45]
  wire [47:0] cluster_59_douta; // @[util.scala 123:45]
  wire  cluster_59_ena; // @[util.scala 123:45]
  wire  cluster_59_wea; // @[util.scala 123:45]
  wire [11:0] cluster_59_addrb; // @[util.scala 123:45]
  wire  cluster_59_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_59_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_59_doutb; // @[util.scala 123:45]
  wire  cluster_59_enb; // @[util.scala 123:45]
  wire  cluster_59_web; // @[util.scala 123:45]
  wire [11:0] cluster_60_addra; // @[util.scala 123:45]
  wire  cluster_60_clka; // @[util.scala 123:45]
  wire [47:0] cluster_60_dina; // @[util.scala 123:45]
  wire [47:0] cluster_60_douta; // @[util.scala 123:45]
  wire  cluster_60_ena; // @[util.scala 123:45]
  wire  cluster_60_wea; // @[util.scala 123:45]
  wire [11:0] cluster_60_addrb; // @[util.scala 123:45]
  wire  cluster_60_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_60_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_60_doutb; // @[util.scala 123:45]
  wire  cluster_60_enb; // @[util.scala 123:45]
  wire  cluster_60_web; // @[util.scala 123:45]
  wire [11:0] cluster_61_addra; // @[util.scala 123:45]
  wire  cluster_61_clka; // @[util.scala 123:45]
  wire [47:0] cluster_61_dina; // @[util.scala 123:45]
  wire [47:0] cluster_61_douta; // @[util.scala 123:45]
  wire  cluster_61_ena; // @[util.scala 123:45]
  wire  cluster_61_wea; // @[util.scala 123:45]
  wire [11:0] cluster_61_addrb; // @[util.scala 123:45]
  wire  cluster_61_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_61_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_61_doutb; // @[util.scala 123:45]
  wire  cluster_61_enb; // @[util.scala 123:45]
  wire  cluster_61_web; // @[util.scala 123:45]
  wire [11:0] cluster_62_addra; // @[util.scala 123:45]
  wire  cluster_62_clka; // @[util.scala 123:45]
  wire [47:0] cluster_62_dina; // @[util.scala 123:45]
  wire [47:0] cluster_62_douta; // @[util.scala 123:45]
  wire  cluster_62_ena; // @[util.scala 123:45]
  wire  cluster_62_wea; // @[util.scala 123:45]
  wire [11:0] cluster_62_addrb; // @[util.scala 123:45]
  wire  cluster_62_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_62_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_62_doutb; // @[util.scala 123:45]
  wire  cluster_62_enb; // @[util.scala 123:45]
  wire  cluster_62_web; // @[util.scala 123:45]
  wire [11:0] cluster_63_addra; // @[util.scala 123:45]
  wire  cluster_63_clka; // @[util.scala 123:45]
  wire [47:0] cluster_63_dina; // @[util.scala 123:45]
  wire [47:0] cluster_63_douta; // @[util.scala 123:45]
  wire  cluster_63_ena; // @[util.scala 123:45]
  wire  cluster_63_wea; // @[util.scala 123:45]
  wire [11:0] cluster_63_addrb; // @[util.scala 123:45]
  wire  cluster_63_clkb; // @[util.scala 123:45]
  wire [47:0] cluster_63_dinb; // @[util.scala 123:45]
  wire [47:0] cluster_63_doutb; // @[util.scala 123:45]
  wire  cluster_63_enb; // @[util.scala 123:45]
  wire  cluster_63_web; // @[util.scala 123:45]
  wire [17:0] _cluster_0_io_web_T = {{12'd0}, io_addrb[17:12]}; // @[util.scala 137:55]
  wire  _cluster_0_io_web_T_1 = 18'h0 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [17:0] _cluster_0_io_wea_T = {{12'd0}, io_addra[17:12]}; // @[util.scala 138:55]
  wire [47:0] doutb_0 = _cluster_0_io_web_T_1 ? cluster_0_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_1_io_web_T_1 = 18'h1 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_1 = _cluster_1_io_web_T_1 ? cluster_1_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_2_io_web_T_1 = 18'h2 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_2 = _cluster_2_io_web_T_1 ? cluster_2_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_3_io_web_T_1 = 18'h3 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_3 = _cluster_3_io_web_T_1 ? cluster_3_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_4_io_web_T_1 = 18'h4 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_4 = _cluster_4_io_web_T_1 ? cluster_4_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_5_io_web_T_1 = 18'h5 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_5 = _cluster_5_io_web_T_1 ? cluster_5_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_6_io_web_T_1 = 18'h6 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_6 = _cluster_6_io_web_T_1 ? cluster_6_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_7_io_web_T_1 = 18'h7 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_7 = _cluster_7_io_web_T_1 ? cluster_7_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_8_io_web_T_1 = 18'h8 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_8 = _cluster_8_io_web_T_1 ? cluster_8_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_9_io_web_T_1 = 18'h9 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_9 = _cluster_9_io_web_T_1 ? cluster_9_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_10_io_web_T_1 = 18'ha == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_10 = _cluster_10_io_web_T_1 ? cluster_10_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_11_io_web_T_1 = 18'hb == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_11 = _cluster_11_io_web_T_1 ? cluster_11_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_12_io_web_T_1 = 18'hc == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_12 = _cluster_12_io_web_T_1 ? cluster_12_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_13_io_web_T_1 = 18'hd == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_13 = _cluster_13_io_web_T_1 ? cluster_13_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_14_io_web_T_1 = 18'he == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_14 = _cluster_14_io_web_T_1 ? cluster_14_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_15_io_web_T_1 = 18'hf == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_15 = _cluster_15_io_web_T_1 ? cluster_15_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_16_io_web_T_1 = 18'h10 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_16 = _cluster_16_io_web_T_1 ? cluster_16_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_17_io_web_T_1 = 18'h11 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_17 = _cluster_17_io_web_T_1 ? cluster_17_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_18_io_web_T_1 = 18'h12 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_18 = _cluster_18_io_web_T_1 ? cluster_18_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_19_io_web_T_1 = 18'h13 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_19 = _cluster_19_io_web_T_1 ? cluster_19_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_20_io_web_T_1 = 18'h14 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_20 = _cluster_20_io_web_T_1 ? cluster_20_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_21_io_web_T_1 = 18'h15 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_21 = _cluster_21_io_web_T_1 ? cluster_21_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_22_io_web_T_1 = 18'h16 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_22 = _cluster_22_io_web_T_1 ? cluster_22_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_23_io_web_T_1 = 18'h17 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_23 = _cluster_23_io_web_T_1 ? cluster_23_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_24_io_web_T_1 = 18'h18 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_24 = _cluster_24_io_web_T_1 ? cluster_24_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_25_io_web_T_1 = 18'h19 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_25 = _cluster_25_io_web_T_1 ? cluster_25_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_26_io_web_T_1 = 18'h1a == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_26 = _cluster_26_io_web_T_1 ? cluster_26_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_27_io_web_T_1 = 18'h1b == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_27 = _cluster_27_io_web_T_1 ? cluster_27_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_28_io_web_T_1 = 18'h1c == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_28 = _cluster_28_io_web_T_1 ? cluster_28_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_29_io_web_T_1 = 18'h1d == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_29 = _cluster_29_io_web_T_1 ? cluster_29_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_30_io_web_T_1 = 18'h1e == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_30 = _cluster_30_io_web_T_1 ? cluster_30_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_31_io_web_T_1 = 18'h1f == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_31 = _cluster_31_io_web_T_1 ? cluster_31_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_32_io_web_T_1 = 18'h20 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_32 = _cluster_32_io_web_T_1 ? cluster_32_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_33_io_web_T_1 = 18'h21 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_33 = _cluster_33_io_web_T_1 ? cluster_33_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_34_io_web_T_1 = 18'h22 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_34 = _cluster_34_io_web_T_1 ? cluster_34_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_35_io_web_T_1 = 18'h23 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_35 = _cluster_35_io_web_T_1 ? cluster_35_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_36_io_web_T_1 = 18'h24 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_36 = _cluster_36_io_web_T_1 ? cluster_36_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_37_io_web_T_1 = 18'h25 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_37 = _cluster_37_io_web_T_1 ? cluster_37_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_38_io_web_T_1 = 18'h26 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_38 = _cluster_38_io_web_T_1 ? cluster_38_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_39_io_web_T_1 = 18'h27 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_39 = _cluster_39_io_web_T_1 ? cluster_39_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_40_io_web_T_1 = 18'h28 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_40 = _cluster_40_io_web_T_1 ? cluster_40_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_41_io_web_T_1 = 18'h29 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_41 = _cluster_41_io_web_T_1 ? cluster_41_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_42_io_web_T_1 = 18'h2a == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_42 = _cluster_42_io_web_T_1 ? cluster_42_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_43_io_web_T_1 = 18'h2b == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_43 = _cluster_43_io_web_T_1 ? cluster_43_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_44_io_web_T_1 = 18'h2c == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_44 = _cluster_44_io_web_T_1 ? cluster_44_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_45_io_web_T_1 = 18'h2d == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_45 = _cluster_45_io_web_T_1 ? cluster_45_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_46_io_web_T_1 = 18'h2e == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_46 = _cluster_46_io_web_T_1 ? cluster_46_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_47_io_web_T_1 = 18'h2f == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_47 = _cluster_47_io_web_T_1 ? cluster_47_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_48_io_web_T_1 = 18'h30 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_48 = _cluster_48_io_web_T_1 ? cluster_48_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_49_io_web_T_1 = 18'h31 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_49 = _cluster_49_io_web_T_1 ? cluster_49_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_50_io_web_T_1 = 18'h32 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_50 = _cluster_50_io_web_T_1 ? cluster_50_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_51_io_web_T_1 = 18'h33 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_51 = _cluster_51_io_web_T_1 ? cluster_51_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_52_io_web_T_1 = 18'h34 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_52 = _cluster_52_io_web_T_1 ? cluster_52_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_53_io_web_T_1 = 18'h35 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_53 = _cluster_53_io_web_T_1 ? cluster_53_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_54_io_web_T_1 = 18'h36 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_54 = _cluster_54_io_web_T_1 ? cluster_54_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_55_io_web_T_1 = 18'h37 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_55 = _cluster_55_io_web_T_1 ? cluster_55_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_56_io_web_T_1 = 18'h38 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_56 = _cluster_56_io_web_T_1 ? cluster_56_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_57_io_web_T_1 = 18'h39 == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_57 = _cluster_57_io_web_T_1 ? cluster_57_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_58_io_web_T_1 = 18'h3a == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_58 = _cluster_58_io_web_T_1 ? cluster_58_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_59_io_web_T_1 = 18'h3b == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_59 = _cluster_59_io_web_T_1 ? cluster_59_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_60_io_web_T_1 = 18'h3c == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_60 = _cluster_60_io_web_T_1 ? cluster_60_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_61_io_web_T_1 = 18'h3d == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_61 = _cluster_61_io_web_T_1 ? cluster_61_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_62_io_web_T_1 = 18'h3e == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_62 = _cluster_62_io_web_T_1 ? cluster_62_doutb : 48'h0; // @[util.scala 139:22]
  wire  _cluster_63_io_web_T_1 = 18'h3f == _cluster_0_io_web_T; // @[util.scala 137:41]
  wire [47:0] doutb_63 = _cluster_63_io_web_T_1 ? cluster_63_doutb : 48'h0; // @[util.scala 139:22]
  wire [47:0] _io_doutb_T = doutb_0 | doutb_1; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_1 = _io_doutb_T | doutb_2; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_2 = _io_doutb_T_1 | doutb_3; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_3 = _io_doutb_T_2 | doutb_4; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_4 = _io_doutb_T_3 | doutb_5; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_5 = _io_doutb_T_4 | doutb_6; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_6 = _io_doutb_T_5 | doutb_7; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_7 = _io_doutb_T_6 | doutb_8; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_8 = _io_doutb_T_7 | doutb_9; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_9 = _io_doutb_T_8 | doutb_10; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_10 = _io_doutb_T_9 | doutb_11; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_11 = _io_doutb_T_10 | doutb_12; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_12 = _io_doutb_T_11 | doutb_13; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_13 = _io_doutb_T_12 | doutb_14; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_14 = _io_doutb_T_13 | doutb_15; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_15 = _io_doutb_T_14 | doutb_16; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_16 = _io_doutb_T_15 | doutb_17; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_17 = _io_doutb_T_16 | doutb_18; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_18 = _io_doutb_T_17 | doutb_19; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_19 = _io_doutb_T_18 | doutb_20; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_20 = _io_doutb_T_19 | doutb_21; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_21 = _io_doutb_T_20 | doutb_22; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_22 = _io_doutb_T_21 | doutb_23; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_23 = _io_doutb_T_22 | doutb_24; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_24 = _io_doutb_T_23 | doutb_25; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_25 = _io_doutb_T_24 | doutb_26; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_26 = _io_doutb_T_25 | doutb_27; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_27 = _io_doutb_T_26 | doutb_28; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_28 = _io_doutb_T_27 | doutb_29; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_29 = _io_doutb_T_28 | doutb_30; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_30 = _io_doutb_T_29 | doutb_31; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_31 = _io_doutb_T_30 | doutb_32; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_32 = _io_doutb_T_31 | doutb_33; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_33 = _io_doutb_T_32 | doutb_34; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_34 = _io_doutb_T_33 | doutb_35; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_35 = _io_doutb_T_34 | doutb_36; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_36 = _io_doutb_T_35 | doutb_37; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_37 = _io_doutb_T_36 | doutb_38; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_38 = _io_doutb_T_37 | doutb_39; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_39 = _io_doutb_T_38 | doutb_40; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_40 = _io_doutb_T_39 | doutb_41; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_41 = _io_doutb_T_40 | doutb_42; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_42 = _io_doutb_T_41 | doutb_43; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_43 = _io_doutb_T_42 | doutb_44; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_44 = _io_doutb_T_43 | doutb_45; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_45 = _io_doutb_T_44 | doutb_46; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_46 = _io_doutb_T_45 | doutb_47; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_47 = _io_doutb_T_46 | doutb_48; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_48 = _io_doutb_T_47 | doutb_49; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_49 = _io_doutb_T_48 | doutb_50; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_50 = _io_doutb_T_49 | doutb_51; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_51 = _io_doutb_T_50 | doutb_52; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_52 = _io_doutb_T_51 | doutb_53; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_53 = _io_doutb_T_52 | doutb_54; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_54 = _io_doutb_T_53 | doutb_55; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_55 = _io_doutb_T_54 | doutb_56; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_56 = _io_doutb_T_55 | doutb_57; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_57 = _io_doutb_T_56 | doutb_58; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_58 = _io_doutb_T_57 | doutb_59; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_59 = _io_doutb_T_58 | doutb_60; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_60 = _io_doutb_T_59 | doutb_61; // @[util.scala 144:29]
  wire [47:0] _io_doutb_T_61 = _io_doutb_T_60 | doutb_62; // @[util.scala 144:29]
  URAM cluster_0 ( // @[util.scala 123:45]
    .addra(cluster_0_addra),
    .clka(cluster_0_clka),
    .dina(cluster_0_dina),
    .douta(cluster_0_douta),
    .ena(cluster_0_ena),
    .wea(cluster_0_wea),
    .addrb(cluster_0_addrb),
    .clkb(cluster_0_clkb),
    .dinb(cluster_0_dinb),
    .doutb(cluster_0_doutb),
    .enb(cluster_0_enb),
    .web(cluster_0_web)
  );
  URAM cluster_1 ( // @[util.scala 123:45]
    .addra(cluster_1_addra),
    .clka(cluster_1_clka),
    .dina(cluster_1_dina),
    .douta(cluster_1_douta),
    .ena(cluster_1_ena),
    .wea(cluster_1_wea),
    .addrb(cluster_1_addrb),
    .clkb(cluster_1_clkb),
    .dinb(cluster_1_dinb),
    .doutb(cluster_1_doutb),
    .enb(cluster_1_enb),
    .web(cluster_1_web)
  );
  URAM cluster_2 ( // @[util.scala 123:45]
    .addra(cluster_2_addra),
    .clka(cluster_2_clka),
    .dina(cluster_2_dina),
    .douta(cluster_2_douta),
    .ena(cluster_2_ena),
    .wea(cluster_2_wea),
    .addrb(cluster_2_addrb),
    .clkb(cluster_2_clkb),
    .dinb(cluster_2_dinb),
    .doutb(cluster_2_doutb),
    .enb(cluster_2_enb),
    .web(cluster_2_web)
  );
  URAM cluster_3 ( // @[util.scala 123:45]
    .addra(cluster_3_addra),
    .clka(cluster_3_clka),
    .dina(cluster_3_dina),
    .douta(cluster_3_douta),
    .ena(cluster_3_ena),
    .wea(cluster_3_wea),
    .addrb(cluster_3_addrb),
    .clkb(cluster_3_clkb),
    .dinb(cluster_3_dinb),
    .doutb(cluster_3_doutb),
    .enb(cluster_3_enb),
    .web(cluster_3_web)
  );
  URAM cluster_4 ( // @[util.scala 123:45]
    .addra(cluster_4_addra),
    .clka(cluster_4_clka),
    .dina(cluster_4_dina),
    .douta(cluster_4_douta),
    .ena(cluster_4_ena),
    .wea(cluster_4_wea),
    .addrb(cluster_4_addrb),
    .clkb(cluster_4_clkb),
    .dinb(cluster_4_dinb),
    .doutb(cluster_4_doutb),
    .enb(cluster_4_enb),
    .web(cluster_4_web)
  );
  URAM cluster_5 ( // @[util.scala 123:45]
    .addra(cluster_5_addra),
    .clka(cluster_5_clka),
    .dina(cluster_5_dina),
    .douta(cluster_5_douta),
    .ena(cluster_5_ena),
    .wea(cluster_5_wea),
    .addrb(cluster_5_addrb),
    .clkb(cluster_5_clkb),
    .dinb(cluster_5_dinb),
    .doutb(cluster_5_doutb),
    .enb(cluster_5_enb),
    .web(cluster_5_web)
  );
  URAM cluster_6 ( // @[util.scala 123:45]
    .addra(cluster_6_addra),
    .clka(cluster_6_clka),
    .dina(cluster_6_dina),
    .douta(cluster_6_douta),
    .ena(cluster_6_ena),
    .wea(cluster_6_wea),
    .addrb(cluster_6_addrb),
    .clkb(cluster_6_clkb),
    .dinb(cluster_6_dinb),
    .doutb(cluster_6_doutb),
    .enb(cluster_6_enb),
    .web(cluster_6_web)
  );
  URAM cluster_7 ( // @[util.scala 123:45]
    .addra(cluster_7_addra),
    .clka(cluster_7_clka),
    .dina(cluster_7_dina),
    .douta(cluster_7_douta),
    .ena(cluster_7_ena),
    .wea(cluster_7_wea),
    .addrb(cluster_7_addrb),
    .clkb(cluster_7_clkb),
    .dinb(cluster_7_dinb),
    .doutb(cluster_7_doutb),
    .enb(cluster_7_enb),
    .web(cluster_7_web)
  );
  URAM cluster_8 ( // @[util.scala 123:45]
    .addra(cluster_8_addra),
    .clka(cluster_8_clka),
    .dina(cluster_8_dina),
    .douta(cluster_8_douta),
    .ena(cluster_8_ena),
    .wea(cluster_8_wea),
    .addrb(cluster_8_addrb),
    .clkb(cluster_8_clkb),
    .dinb(cluster_8_dinb),
    .doutb(cluster_8_doutb),
    .enb(cluster_8_enb),
    .web(cluster_8_web)
  );
  URAM cluster_9 ( // @[util.scala 123:45]
    .addra(cluster_9_addra),
    .clka(cluster_9_clka),
    .dina(cluster_9_dina),
    .douta(cluster_9_douta),
    .ena(cluster_9_ena),
    .wea(cluster_9_wea),
    .addrb(cluster_9_addrb),
    .clkb(cluster_9_clkb),
    .dinb(cluster_9_dinb),
    .doutb(cluster_9_doutb),
    .enb(cluster_9_enb),
    .web(cluster_9_web)
  );
  URAM cluster_10 ( // @[util.scala 123:45]
    .addra(cluster_10_addra),
    .clka(cluster_10_clka),
    .dina(cluster_10_dina),
    .douta(cluster_10_douta),
    .ena(cluster_10_ena),
    .wea(cluster_10_wea),
    .addrb(cluster_10_addrb),
    .clkb(cluster_10_clkb),
    .dinb(cluster_10_dinb),
    .doutb(cluster_10_doutb),
    .enb(cluster_10_enb),
    .web(cluster_10_web)
  );
  URAM cluster_11 ( // @[util.scala 123:45]
    .addra(cluster_11_addra),
    .clka(cluster_11_clka),
    .dina(cluster_11_dina),
    .douta(cluster_11_douta),
    .ena(cluster_11_ena),
    .wea(cluster_11_wea),
    .addrb(cluster_11_addrb),
    .clkb(cluster_11_clkb),
    .dinb(cluster_11_dinb),
    .doutb(cluster_11_doutb),
    .enb(cluster_11_enb),
    .web(cluster_11_web)
  );
  URAM cluster_12 ( // @[util.scala 123:45]
    .addra(cluster_12_addra),
    .clka(cluster_12_clka),
    .dina(cluster_12_dina),
    .douta(cluster_12_douta),
    .ena(cluster_12_ena),
    .wea(cluster_12_wea),
    .addrb(cluster_12_addrb),
    .clkb(cluster_12_clkb),
    .dinb(cluster_12_dinb),
    .doutb(cluster_12_doutb),
    .enb(cluster_12_enb),
    .web(cluster_12_web)
  );
  URAM cluster_13 ( // @[util.scala 123:45]
    .addra(cluster_13_addra),
    .clka(cluster_13_clka),
    .dina(cluster_13_dina),
    .douta(cluster_13_douta),
    .ena(cluster_13_ena),
    .wea(cluster_13_wea),
    .addrb(cluster_13_addrb),
    .clkb(cluster_13_clkb),
    .dinb(cluster_13_dinb),
    .doutb(cluster_13_doutb),
    .enb(cluster_13_enb),
    .web(cluster_13_web)
  );
  URAM cluster_14 ( // @[util.scala 123:45]
    .addra(cluster_14_addra),
    .clka(cluster_14_clka),
    .dina(cluster_14_dina),
    .douta(cluster_14_douta),
    .ena(cluster_14_ena),
    .wea(cluster_14_wea),
    .addrb(cluster_14_addrb),
    .clkb(cluster_14_clkb),
    .dinb(cluster_14_dinb),
    .doutb(cluster_14_doutb),
    .enb(cluster_14_enb),
    .web(cluster_14_web)
  );
  URAM cluster_15 ( // @[util.scala 123:45]
    .addra(cluster_15_addra),
    .clka(cluster_15_clka),
    .dina(cluster_15_dina),
    .douta(cluster_15_douta),
    .ena(cluster_15_ena),
    .wea(cluster_15_wea),
    .addrb(cluster_15_addrb),
    .clkb(cluster_15_clkb),
    .dinb(cluster_15_dinb),
    .doutb(cluster_15_doutb),
    .enb(cluster_15_enb),
    .web(cluster_15_web)
  );
  URAM cluster_16 ( // @[util.scala 123:45]
    .addra(cluster_16_addra),
    .clka(cluster_16_clka),
    .dina(cluster_16_dina),
    .douta(cluster_16_douta),
    .ena(cluster_16_ena),
    .wea(cluster_16_wea),
    .addrb(cluster_16_addrb),
    .clkb(cluster_16_clkb),
    .dinb(cluster_16_dinb),
    .doutb(cluster_16_doutb),
    .enb(cluster_16_enb),
    .web(cluster_16_web)
  );
  URAM cluster_17 ( // @[util.scala 123:45]
    .addra(cluster_17_addra),
    .clka(cluster_17_clka),
    .dina(cluster_17_dina),
    .douta(cluster_17_douta),
    .ena(cluster_17_ena),
    .wea(cluster_17_wea),
    .addrb(cluster_17_addrb),
    .clkb(cluster_17_clkb),
    .dinb(cluster_17_dinb),
    .doutb(cluster_17_doutb),
    .enb(cluster_17_enb),
    .web(cluster_17_web)
  );
  URAM cluster_18 ( // @[util.scala 123:45]
    .addra(cluster_18_addra),
    .clka(cluster_18_clka),
    .dina(cluster_18_dina),
    .douta(cluster_18_douta),
    .ena(cluster_18_ena),
    .wea(cluster_18_wea),
    .addrb(cluster_18_addrb),
    .clkb(cluster_18_clkb),
    .dinb(cluster_18_dinb),
    .doutb(cluster_18_doutb),
    .enb(cluster_18_enb),
    .web(cluster_18_web)
  );
  URAM cluster_19 ( // @[util.scala 123:45]
    .addra(cluster_19_addra),
    .clka(cluster_19_clka),
    .dina(cluster_19_dina),
    .douta(cluster_19_douta),
    .ena(cluster_19_ena),
    .wea(cluster_19_wea),
    .addrb(cluster_19_addrb),
    .clkb(cluster_19_clkb),
    .dinb(cluster_19_dinb),
    .doutb(cluster_19_doutb),
    .enb(cluster_19_enb),
    .web(cluster_19_web)
  );
  URAM cluster_20 ( // @[util.scala 123:45]
    .addra(cluster_20_addra),
    .clka(cluster_20_clka),
    .dina(cluster_20_dina),
    .douta(cluster_20_douta),
    .ena(cluster_20_ena),
    .wea(cluster_20_wea),
    .addrb(cluster_20_addrb),
    .clkb(cluster_20_clkb),
    .dinb(cluster_20_dinb),
    .doutb(cluster_20_doutb),
    .enb(cluster_20_enb),
    .web(cluster_20_web)
  );
  URAM cluster_21 ( // @[util.scala 123:45]
    .addra(cluster_21_addra),
    .clka(cluster_21_clka),
    .dina(cluster_21_dina),
    .douta(cluster_21_douta),
    .ena(cluster_21_ena),
    .wea(cluster_21_wea),
    .addrb(cluster_21_addrb),
    .clkb(cluster_21_clkb),
    .dinb(cluster_21_dinb),
    .doutb(cluster_21_doutb),
    .enb(cluster_21_enb),
    .web(cluster_21_web)
  );
  URAM cluster_22 ( // @[util.scala 123:45]
    .addra(cluster_22_addra),
    .clka(cluster_22_clka),
    .dina(cluster_22_dina),
    .douta(cluster_22_douta),
    .ena(cluster_22_ena),
    .wea(cluster_22_wea),
    .addrb(cluster_22_addrb),
    .clkb(cluster_22_clkb),
    .dinb(cluster_22_dinb),
    .doutb(cluster_22_doutb),
    .enb(cluster_22_enb),
    .web(cluster_22_web)
  );
  URAM cluster_23 ( // @[util.scala 123:45]
    .addra(cluster_23_addra),
    .clka(cluster_23_clka),
    .dina(cluster_23_dina),
    .douta(cluster_23_douta),
    .ena(cluster_23_ena),
    .wea(cluster_23_wea),
    .addrb(cluster_23_addrb),
    .clkb(cluster_23_clkb),
    .dinb(cluster_23_dinb),
    .doutb(cluster_23_doutb),
    .enb(cluster_23_enb),
    .web(cluster_23_web)
  );
  URAM cluster_24 ( // @[util.scala 123:45]
    .addra(cluster_24_addra),
    .clka(cluster_24_clka),
    .dina(cluster_24_dina),
    .douta(cluster_24_douta),
    .ena(cluster_24_ena),
    .wea(cluster_24_wea),
    .addrb(cluster_24_addrb),
    .clkb(cluster_24_clkb),
    .dinb(cluster_24_dinb),
    .doutb(cluster_24_doutb),
    .enb(cluster_24_enb),
    .web(cluster_24_web)
  );
  URAM cluster_25 ( // @[util.scala 123:45]
    .addra(cluster_25_addra),
    .clka(cluster_25_clka),
    .dina(cluster_25_dina),
    .douta(cluster_25_douta),
    .ena(cluster_25_ena),
    .wea(cluster_25_wea),
    .addrb(cluster_25_addrb),
    .clkb(cluster_25_clkb),
    .dinb(cluster_25_dinb),
    .doutb(cluster_25_doutb),
    .enb(cluster_25_enb),
    .web(cluster_25_web)
  );
  URAM cluster_26 ( // @[util.scala 123:45]
    .addra(cluster_26_addra),
    .clka(cluster_26_clka),
    .dina(cluster_26_dina),
    .douta(cluster_26_douta),
    .ena(cluster_26_ena),
    .wea(cluster_26_wea),
    .addrb(cluster_26_addrb),
    .clkb(cluster_26_clkb),
    .dinb(cluster_26_dinb),
    .doutb(cluster_26_doutb),
    .enb(cluster_26_enb),
    .web(cluster_26_web)
  );
  URAM cluster_27 ( // @[util.scala 123:45]
    .addra(cluster_27_addra),
    .clka(cluster_27_clka),
    .dina(cluster_27_dina),
    .douta(cluster_27_douta),
    .ena(cluster_27_ena),
    .wea(cluster_27_wea),
    .addrb(cluster_27_addrb),
    .clkb(cluster_27_clkb),
    .dinb(cluster_27_dinb),
    .doutb(cluster_27_doutb),
    .enb(cluster_27_enb),
    .web(cluster_27_web)
  );
  URAM cluster_28 ( // @[util.scala 123:45]
    .addra(cluster_28_addra),
    .clka(cluster_28_clka),
    .dina(cluster_28_dina),
    .douta(cluster_28_douta),
    .ena(cluster_28_ena),
    .wea(cluster_28_wea),
    .addrb(cluster_28_addrb),
    .clkb(cluster_28_clkb),
    .dinb(cluster_28_dinb),
    .doutb(cluster_28_doutb),
    .enb(cluster_28_enb),
    .web(cluster_28_web)
  );
  URAM cluster_29 ( // @[util.scala 123:45]
    .addra(cluster_29_addra),
    .clka(cluster_29_clka),
    .dina(cluster_29_dina),
    .douta(cluster_29_douta),
    .ena(cluster_29_ena),
    .wea(cluster_29_wea),
    .addrb(cluster_29_addrb),
    .clkb(cluster_29_clkb),
    .dinb(cluster_29_dinb),
    .doutb(cluster_29_doutb),
    .enb(cluster_29_enb),
    .web(cluster_29_web)
  );
  URAM cluster_30 ( // @[util.scala 123:45]
    .addra(cluster_30_addra),
    .clka(cluster_30_clka),
    .dina(cluster_30_dina),
    .douta(cluster_30_douta),
    .ena(cluster_30_ena),
    .wea(cluster_30_wea),
    .addrb(cluster_30_addrb),
    .clkb(cluster_30_clkb),
    .dinb(cluster_30_dinb),
    .doutb(cluster_30_doutb),
    .enb(cluster_30_enb),
    .web(cluster_30_web)
  );
  URAM cluster_31 ( // @[util.scala 123:45]
    .addra(cluster_31_addra),
    .clka(cluster_31_clka),
    .dina(cluster_31_dina),
    .douta(cluster_31_douta),
    .ena(cluster_31_ena),
    .wea(cluster_31_wea),
    .addrb(cluster_31_addrb),
    .clkb(cluster_31_clkb),
    .dinb(cluster_31_dinb),
    .doutb(cluster_31_doutb),
    .enb(cluster_31_enb),
    .web(cluster_31_web)
  );
  URAM cluster_32 ( // @[util.scala 123:45]
    .addra(cluster_32_addra),
    .clka(cluster_32_clka),
    .dina(cluster_32_dina),
    .douta(cluster_32_douta),
    .ena(cluster_32_ena),
    .wea(cluster_32_wea),
    .addrb(cluster_32_addrb),
    .clkb(cluster_32_clkb),
    .dinb(cluster_32_dinb),
    .doutb(cluster_32_doutb),
    .enb(cluster_32_enb),
    .web(cluster_32_web)
  );
  URAM cluster_33 ( // @[util.scala 123:45]
    .addra(cluster_33_addra),
    .clka(cluster_33_clka),
    .dina(cluster_33_dina),
    .douta(cluster_33_douta),
    .ena(cluster_33_ena),
    .wea(cluster_33_wea),
    .addrb(cluster_33_addrb),
    .clkb(cluster_33_clkb),
    .dinb(cluster_33_dinb),
    .doutb(cluster_33_doutb),
    .enb(cluster_33_enb),
    .web(cluster_33_web)
  );
  URAM cluster_34 ( // @[util.scala 123:45]
    .addra(cluster_34_addra),
    .clka(cluster_34_clka),
    .dina(cluster_34_dina),
    .douta(cluster_34_douta),
    .ena(cluster_34_ena),
    .wea(cluster_34_wea),
    .addrb(cluster_34_addrb),
    .clkb(cluster_34_clkb),
    .dinb(cluster_34_dinb),
    .doutb(cluster_34_doutb),
    .enb(cluster_34_enb),
    .web(cluster_34_web)
  );
  URAM cluster_35 ( // @[util.scala 123:45]
    .addra(cluster_35_addra),
    .clka(cluster_35_clka),
    .dina(cluster_35_dina),
    .douta(cluster_35_douta),
    .ena(cluster_35_ena),
    .wea(cluster_35_wea),
    .addrb(cluster_35_addrb),
    .clkb(cluster_35_clkb),
    .dinb(cluster_35_dinb),
    .doutb(cluster_35_doutb),
    .enb(cluster_35_enb),
    .web(cluster_35_web)
  );
  URAM cluster_36 ( // @[util.scala 123:45]
    .addra(cluster_36_addra),
    .clka(cluster_36_clka),
    .dina(cluster_36_dina),
    .douta(cluster_36_douta),
    .ena(cluster_36_ena),
    .wea(cluster_36_wea),
    .addrb(cluster_36_addrb),
    .clkb(cluster_36_clkb),
    .dinb(cluster_36_dinb),
    .doutb(cluster_36_doutb),
    .enb(cluster_36_enb),
    .web(cluster_36_web)
  );
  URAM cluster_37 ( // @[util.scala 123:45]
    .addra(cluster_37_addra),
    .clka(cluster_37_clka),
    .dina(cluster_37_dina),
    .douta(cluster_37_douta),
    .ena(cluster_37_ena),
    .wea(cluster_37_wea),
    .addrb(cluster_37_addrb),
    .clkb(cluster_37_clkb),
    .dinb(cluster_37_dinb),
    .doutb(cluster_37_doutb),
    .enb(cluster_37_enb),
    .web(cluster_37_web)
  );
  URAM cluster_38 ( // @[util.scala 123:45]
    .addra(cluster_38_addra),
    .clka(cluster_38_clka),
    .dina(cluster_38_dina),
    .douta(cluster_38_douta),
    .ena(cluster_38_ena),
    .wea(cluster_38_wea),
    .addrb(cluster_38_addrb),
    .clkb(cluster_38_clkb),
    .dinb(cluster_38_dinb),
    .doutb(cluster_38_doutb),
    .enb(cluster_38_enb),
    .web(cluster_38_web)
  );
  URAM cluster_39 ( // @[util.scala 123:45]
    .addra(cluster_39_addra),
    .clka(cluster_39_clka),
    .dina(cluster_39_dina),
    .douta(cluster_39_douta),
    .ena(cluster_39_ena),
    .wea(cluster_39_wea),
    .addrb(cluster_39_addrb),
    .clkb(cluster_39_clkb),
    .dinb(cluster_39_dinb),
    .doutb(cluster_39_doutb),
    .enb(cluster_39_enb),
    .web(cluster_39_web)
  );
  URAM cluster_40 ( // @[util.scala 123:45]
    .addra(cluster_40_addra),
    .clka(cluster_40_clka),
    .dina(cluster_40_dina),
    .douta(cluster_40_douta),
    .ena(cluster_40_ena),
    .wea(cluster_40_wea),
    .addrb(cluster_40_addrb),
    .clkb(cluster_40_clkb),
    .dinb(cluster_40_dinb),
    .doutb(cluster_40_doutb),
    .enb(cluster_40_enb),
    .web(cluster_40_web)
  );
  URAM cluster_41 ( // @[util.scala 123:45]
    .addra(cluster_41_addra),
    .clka(cluster_41_clka),
    .dina(cluster_41_dina),
    .douta(cluster_41_douta),
    .ena(cluster_41_ena),
    .wea(cluster_41_wea),
    .addrb(cluster_41_addrb),
    .clkb(cluster_41_clkb),
    .dinb(cluster_41_dinb),
    .doutb(cluster_41_doutb),
    .enb(cluster_41_enb),
    .web(cluster_41_web)
  );
  URAM cluster_42 ( // @[util.scala 123:45]
    .addra(cluster_42_addra),
    .clka(cluster_42_clka),
    .dina(cluster_42_dina),
    .douta(cluster_42_douta),
    .ena(cluster_42_ena),
    .wea(cluster_42_wea),
    .addrb(cluster_42_addrb),
    .clkb(cluster_42_clkb),
    .dinb(cluster_42_dinb),
    .doutb(cluster_42_doutb),
    .enb(cluster_42_enb),
    .web(cluster_42_web)
  );
  URAM cluster_43 ( // @[util.scala 123:45]
    .addra(cluster_43_addra),
    .clka(cluster_43_clka),
    .dina(cluster_43_dina),
    .douta(cluster_43_douta),
    .ena(cluster_43_ena),
    .wea(cluster_43_wea),
    .addrb(cluster_43_addrb),
    .clkb(cluster_43_clkb),
    .dinb(cluster_43_dinb),
    .doutb(cluster_43_doutb),
    .enb(cluster_43_enb),
    .web(cluster_43_web)
  );
  URAM cluster_44 ( // @[util.scala 123:45]
    .addra(cluster_44_addra),
    .clka(cluster_44_clka),
    .dina(cluster_44_dina),
    .douta(cluster_44_douta),
    .ena(cluster_44_ena),
    .wea(cluster_44_wea),
    .addrb(cluster_44_addrb),
    .clkb(cluster_44_clkb),
    .dinb(cluster_44_dinb),
    .doutb(cluster_44_doutb),
    .enb(cluster_44_enb),
    .web(cluster_44_web)
  );
  URAM cluster_45 ( // @[util.scala 123:45]
    .addra(cluster_45_addra),
    .clka(cluster_45_clka),
    .dina(cluster_45_dina),
    .douta(cluster_45_douta),
    .ena(cluster_45_ena),
    .wea(cluster_45_wea),
    .addrb(cluster_45_addrb),
    .clkb(cluster_45_clkb),
    .dinb(cluster_45_dinb),
    .doutb(cluster_45_doutb),
    .enb(cluster_45_enb),
    .web(cluster_45_web)
  );
  URAM cluster_46 ( // @[util.scala 123:45]
    .addra(cluster_46_addra),
    .clka(cluster_46_clka),
    .dina(cluster_46_dina),
    .douta(cluster_46_douta),
    .ena(cluster_46_ena),
    .wea(cluster_46_wea),
    .addrb(cluster_46_addrb),
    .clkb(cluster_46_clkb),
    .dinb(cluster_46_dinb),
    .doutb(cluster_46_doutb),
    .enb(cluster_46_enb),
    .web(cluster_46_web)
  );
  URAM cluster_47 ( // @[util.scala 123:45]
    .addra(cluster_47_addra),
    .clka(cluster_47_clka),
    .dina(cluster_47_dina),
    .douta(cluster_47_douta),
    .ena(cluster_47_ena),
    .wea(cluster_47_wea),
    .addrb(cluster_47_addrb),
    .clkb(cluster_47_clkb),
    .dinb(cluster_47_dinb),
    .doutb(cluster_47_doutb),
    .enb(cluster_47_enb),
    .web(cluster_47_web)
  );
  URAM cluster_48 ( // @[util.scala 123:45]
    .addra(cluster_48_addra),
    .clka(cluster_48_clka),
    .dina(cluster_48_dina),
    .douta(cluster_48_douta),
    .ena(cluster_48_ena),
    .wea(cluster_48_wea),
    .addrb(cluster_48_addrb),
    .clkb(cluster_48_clkb),
    .dinb(cluster_48_dinb),
    .doutb(cluster_48_doutb),
    .enb(cluster_48_enb),
    .web(cluster_48_web)
  );
  URAM cluster_49 ( // @[util.scala 123:45]
    .addra(cluster_49_addra),
    .clka(cluster_49_clka),
    .dina(cluster_49_dina),
    .douta(cluster_49_douta),
    .ena(cluster_49_ena),
    .wea(cluster_49_wea),
    .addrb(cluster_49_addrb),
    .clkb(cluster_49_clkb),
    .dinb(cluster_49_dinb),
    .doutb(cluster_49_doutb),
    .enb(cluster_49_enb),
    .web(cluster_49_web)
  );
  URAM cluster_50 ( // @[util.scala 123:45]
    .addra(cluster_50_addra),
    .clka(cluster_50_clka),
    .dina(cluster_50_dina),
    .douta(cluster_50_douta),
    .ena(cluster_50_ena),
    .wea(cluster_50_wea),
    .addrb(cluster_50_addrb),
    .clkb(cluster_50_clkb),
    .dinb(cluster_50_dinb),
    .doutb(cluster_50_doutb),
    .enb(cluster_50_enb),
    .web(cluster_50_web)
  );
  URAM cluster_51 ( // @[util.scala 123:45]
    .addra(cluster_51_addra),
    .clka(cluster_51_clka),
    .dina(cluster_51_dina),
    .douta(cluster_51_douta),
    .ena(cluster_51_ena),
    .wea(cluster_51_wea),
    .addrb(cluster_51_addrb),
    .clkb(cluster_51_clkb),
    .dinb(cluster_51_dinb),
    .doutb(cluster_51_doutb),
    .enb(cluster_51_enb),
    .web(cluster_51_web)
  );
  URAM cluster_52 ( // @[util.scala 123:45]
    .addra(cluster_52_addra),
    .clka(cluster_52_clka),
    .dina(cluster_52_dina),
    .douta(cluster_52_douta),
    .ena(cluster_52_ena),
    .wea(cluster_52_wea),
    .addrb(cluster_52_addrb),
    .clkb(cluster_52_clkb),
    .dinb(cluster_52_dinb),
    .doutb(cluster_52_doutb),
    .enb(cluster_52_enb),
    .web(cluster_52_web)
  );
  URAM cluster_53 ( // @[util.scala 123:45]
    .addra(cluster_53_addra),
    .clka(cluster_53_clka),
    .dina(cluster_53_dina),
    .douta(cluster_53_douta),
    .ena(cluster_53_ena),
    .wea(cluster_53_wea),
    .addrb(cluster_53_addrb),
    .clkb(cluster_53_clkb),
    .dinb(cluster_53_dinb),
    .doutb(cluster_53_doutb),
    .enb(cluster_53_enb),
    .web(cluster_53_web)
  );
  URAM cluster_54 ( // @[util.scala 123:45]
    .addra(cluster_54_addra),
    .clka(cluster_54_clka),
    .dina(cluster_54_dina),
    .douta(cluster_54_douta),
    .ena(cluster_54_ena),
    .wea(cluster_54_wea),
    .addrb(cluster_54_addrb),
    .clkb(cluster_54_clkb),
    .dinb(cluster_54_dinb),
    .doutb(cluster_54_doutb),
    .enb(cluster_54_enb),
    .web(cluster_54_web)
  );
  URAM cluster_55 ( // @[util.scala 123:45]
    .addra(cluster_55_addra),
    .clka(cluster_55_clka),
    .dina(cluster_55_dina),
    .douta(cluster_55_douta),
    .ena(cluster_55_ena),
    .wea(cluster_55_wea),
    .addrb(cluster_55_addrb),
    .clkb(cluster_55_clkb),
    .dinb(cluster_55_dinb),
    .doutb(cluster_55_doutb),
    .enb(cluster_55_enb),
    .web(cluster_55_web)
  );
  URAM cluster_56 ( // @[util.scala 123:45]
    .addra(cluster_56_addra),
    .clka(cluster_56_clka),
    .dina(cluster_56_dina),
    .douta(cluster_56_douta),
    .ena(cluster_56_ena),
    .wea(cluster_56_wea),
    .addrb(cluster_56_addrb),
    .clkb(cluster_56_clkb),
    .dinb(cluster_56_dinb),
    .doutb(cluster_56_doutb),
    .enb(cluster_56_enb),
    .web(cluster_56_web)
  );
  URAM cluster_57 ( // @[util.scala 123:45]
    .addra(cluster_57_addra),
    .clka(cluster_57_clka),
    .dina(cluster_57_dina),
    .douta(cluster_57_douta),
    .ena(cluster_57_ena),
    .wea(cluster_57_wea),
    .addrb(cluster_57_addrb),
    .clkb(cluster_57_clkb),
    .dinb(cluster_57_dinb),
    .doutb(cluster_57_doutb),
    .enb(cluster_57_enb),
    .web(cluster_57_web)
  );
  URAM cluster_58 ( // @[util.scala 123:45]
    .addra(cluster_58_addra),
    .clka(cluster_58_clka),
    .dina(cluster_58_dina),
    .douta(cluster_58_douta),
    .ena(cluster_58_ena),
    .wea(cluster_58_wea),
    .addrb(cluster_58_addrb),
    .clkb(cluster_58_clkb),
    .dinb(cluster_58_dinb),
    .doutb(cluster_58_doutb),
    .enb(cluster_58_enb),
    .web(cluster_58_web)
  );
  URAM cluster_59 ( // @[util.scala 123:45]
    .addra(cluster_59_addra),
    .clka(cluster_59_clka),
    .dina(cluster_59_dina),
    .douta(cluster_59_douta),
    .ena(cluster_59_ena),
    .wea(cluster_59_wea),
    .addrb(cluster_59_addrb),
    .clkb(cluster_59_clkb),
    .dinb(cluster_59_dinb),
    .doutb(cluster_59_doutb),
    .enb(cluster_59_enb),
    .web(cluster_59_web)
  );
  URAM cluster_60 ( // @[util.scala 123:45]
    .addra(cluster_60_addra),
    .clka(cluster_60_clka),
    .dina(cluster_60_dina),
    .douta(cluster_60_douta),
    .ena(cluster_60_ena),
    .wea(cluster_60_wea),
    .addrb(cluster_60_addrb),
    .clkb(cluster_60_clkb),
    .dinb(cluster_60_dinb),
    .doutb(cluster_60_doutb),
    .enb(cluster_60_enb),
    .web(cluster_60_web)
  );
  URAM cluster_61 ( // @[util.scala 123:45]
    .addra(cluster_61_addra),
    .clka(cluster_61_clka),
    .dina(cluster_61_dina),
    .douta(cluster_61_douta),
    .ena(cluster_61_ena),
    .wea(cluster_61_wea),
    .addrb(cluster_61_addrb),
    .clkb(cluster_61_clkb),
    .dinb(cluster_61_dinb),
    .doutb(cluster_61_doutb),
    .enb(cluster_61_enb),
    .web(cluster_61_web)
  );
  URAM cluster_62 ( // @[util.scala 123:45]
    .addra(cluster_62_addra),
    .clka(cluster_62_clka),
    .dina(cluster_62_dina),
    .douta(cluster_62_douta),
    .ena(cluster_62_ena),
    .wea(cluster_62_wea),
    .addrb(cluster_62_addrb),
    .clkb(cluster_62_clkb),
    .dinb(cluster_62_dinb),
    .doutb(cluster_62_doutb),
    .enb(cluster_62_enb),
    .web(cluster_62_web)
  );
  URAM cluster_63 ( // @[util.scala 123:45]
    .addra(cluster_63_addra),
    .clka(cluster_63_clka),
    .dina(cluster_63_dina),
    .douta(cluster_63_douta),
    .ena(cluster_63_ena),
    .wea(cluster_63_wea),
    .addrb(cluster_63_addrb),
    .clkb(cluster_63_clkb),
    .dinb(cluster_63_dinb),
    .doutb(cluster_63_doutb),
    .enb(cluster_63_enb),
    .web(cluster_63_web)
  );
  assign io_doutb = _io_doutb_T_61 | doutb_63; // @[util.scala 144:29]
  assign cluster_0_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_0_clka = io_clka; // @[util.scala 130:17]
  assign cluster_0_dina = io_dina; // @[util.scala 134:17]
  assign cluster_0_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_0_wea = io_wea & 18'h0 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_0_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_0_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_0_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_0_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_0_web = 1'h0; // @[util.scala 137:26]
  assign cluster_1_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_1_clka = io_clka; // @[util.scala 130:17]
  assign cluster_1_dina = io_dina; // @[util.scala 134:17]
  assign cluster_1_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_1_wea = io_wea & 18'h1 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_1_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_1_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_1_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_1_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_1_web = 1'h0; // @[util.scala 137:26]
  assign cluster_2_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_2_clka = io_clka; // @[util.scala 130:17]
  assign cluster_2_dina = io_dina; // @[util.scala 134:17]
  assign cluster_2_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_2_wea = io_wea & 18'h2 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_2_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_2_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_2_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_2_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_2_web = 1'h0; // @[util.scala 137:26]
  assign cluster_3_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_3_clka = io_clka; // @[util.scala 130:17]
  assign cluster_3_dina = io_dina; // @[util.scala 134:17]
  assign cluster_3_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_3_wea = io_wea & 18'h3 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_3_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_3_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_3_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_3_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_3_web = 1'h0; // @[util.scala 137:26]
  assign cluster_4_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_4_clka = io_clka; // @[util.scala 130:17]
  assign cluster_4_dina = io_dina; // @[util.scala 134:17]
  assign cluster_4_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_4_wea = io_wea & 18'h4 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_4_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_4_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_4_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_4_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_4_web = 1'h0; // @[util.scala 137:26]
  assign cluster_5_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_5_clka = io_clka; // @[util.scala 130:17]
  assign cluster_5_dina = io_dina; // @[util.scala 134:17]
  assign cluster_5_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_5_wea = io_wea & 18'h5 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_5_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_5_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_5_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_5_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_5_web = 1'h0; // @[util.scala 137:26]
  assign cluster_6_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_6_clka = io_clka; // @[util.scala 130:17]
  assign cluster_6_dina = io_dina; // @[util.scala 134:17]
  assign cluster_6_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_6_wea = io_wea & 18'h6 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_6_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_6_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_6_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_6_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_6_web = 1'h0; // @[util.scala 137:26]
  assign cluster_7_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_7_clka = io_clka; // @[util.scala 130:17]
  assign cluster_7_dina = io_dina; // @[util.scala 134:17]
  assign cluster_7_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_7_wea = io_wea & 18'h7 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_7_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_7_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_7_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_7_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_7_web = 1'h0; // @[util.scala 137:26]
  assign cluster_8_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_8_clka = io_clka; // @[util.scala 130:17]
  assign cluster_8_dina = io_dina; // @[util.scala 134:17]
  assign cluster_8_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_8_wea = io_wea & 18'h8 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_8_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_8_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_8_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_8_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_8_web = 1'h0; // @[util.scala 137:26]
  assign cluster_9_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_9_clka = io_clka; // @[util.scala 130:17]
  assign cluster_9_dina = io_dina; // @[util.scala 134:17]
  assign cluster_9_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_9_wea = io_wea & 18'h9 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_9_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_9_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_9_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_9_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_9_web = 1'h0; // @[util.scala 137:26]
  assign cluster_10_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_10_clka = io_clka; // @[util.scala 130:17]
  assign cluster_10_dina = io_dina; // @[util.scala 134:17]
  assign cluster_10_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_10_wea = io_wea & 18'ha == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_10_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_10_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_10_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_10_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_10_web = 1'h0; // @[util.scala 137:26]
  assign cluster_11_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_11_clka = io_clka; // @[util.scala 130:17]
  assign cluster_11_dina = io_dina; // @[util.scala 134:17]
  assign cluster_11_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_11_wea = io_wea & 18'hb == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_11_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_11_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_11_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_11_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_11_web = 1'h0; // @[util.scala 137:26]
  assign cluster_12_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_12_clka = io_clka; // @[util.scala 130:17]
  assign cluster_12_dina = io_dina; // @[util.scala 134:17]
  assign cluster_12_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_12_wea = io_wea & 18'hc == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_12_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_12_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_12_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_12_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_12_web = 1'h0; // @[util.scala 137:26]
  assign cluster_13_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_13_clka = io_clka; // @[util.scala 130:17]
  assign cluster_13_dina = io_dina; // @[util.scala 134:17]
  assign cluster_13_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_13_wea = io_wea & 18'hd == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_13_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_13_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_13_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_13_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_13_web = 1'h0; // @[util.scala 137:26]
  assign cluster_14_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_14_clka = io_clka; // @[util.scala 130:17]
  assign cluster_14_dina = io_dina; // @[util.scala 134:17]
  assign cluster_14_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_14_wea = io_wea & 18'he == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_14_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_14_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_14_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_14_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_14_web = 1'h0; // @[util.scala 137:26]
  assign cluster_15_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_15_clka = io_clka; // @[util.scala 130:17]
  assign cluster_15_dina = io_dina; // @[util.scala 134:17]
  assign cluster_15_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_15_wea = io_wea & 18'hf == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_15_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_15_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_15_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_15_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_15_web = 1'h0; // @[util.scala 137:26]
  assign cluster_16_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_16_clka = io_clka; // @[util.scala 130:17]
  assign cluster_16_dina = io_dina; // @[util.scala 134:17]
  assign cluster_16_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_16_wea = io_wea & 18'h10 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_16_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_16_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_16_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_16_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_16_web = 1'h0; // @[util.scala 137:26]
  assign cluster_17_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_17_clka = io_clka; // @[util.scala 130:17]
  assign cluster_17_dina = io_dina; // @[util.scala 134:17]
  assign cluster_17_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_17_wea = io_wea & 18'h11 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_17_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_17_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_17_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_17_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_17_web = 1'h0; // @[util.scala 137:26]
  assign cluster_18_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_18_clka = io_clka; // @[util.scala 130:17]
  assign cluster_18_dina = io_dina; // @[util.scala 134:17]
  assign cluster_18_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_18_wea = io_wea & 18'h12 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_18_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_18_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_18_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_18_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_18_web = 1'h0; // @[util.scala 137:26]
  assign cluster_19_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_19_clka = io_clka; // @[util.scala 130:17]
  assign cluster_19_dina = io_dina; // @[util.scala 134:17]
  assign cluster_19_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_19_wea = io_wea & 18'h13 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_19_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_19_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_19_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_19_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_19_web = 1'h0; // @[util.scala 137:26]
  assign cluster_20_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_20_clka = io_clka; // @[util.scala 130:17]
  assign cluster_20_dina = io_dina; // @[util.scala 134:17]
  assign cluster_20_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_20_wea = io_wea & 18'h14 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_20_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_20_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_20_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_20_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_20_web = 1'h0; // @[util.scala 137:26]
  assign cluster_21_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_21_clka = io_clka; // @[util.scala 130:17]
  assign cluster_21_dina = io_dina; // @[util.scala 134:17]
  assign cluster_21_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_21_wea = io_wea & 18'h15 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_21_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_21_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_21_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_21_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_21_web = 1'h0; // @[util.scala 137:26]
  assign cluster_22_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_22_clka = io_clka; // @[util.scala 130:17]
  assign cluster_22_dina = io_dina; // @[util.scala 134:17]
  assign cluster_22_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_22_wea = io_wea & 18'h16 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_22_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_22_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_22_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_22_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_22_web = 1'h0; // @[util.scala 137:26]
  assign cluster_23_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_23_clka = io_clka; // @[util.scala 130:17]
  assign cluster_23_dina = io_dina; // @[util.scala 134:17]
  assign cluster_23_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_23_wea = io_wea & 18'h17 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_23_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_23_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_23_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_23_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_23_web = 1'h0; // @[util.scala 137:26]
  assign cluster_24_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_24_clka = io_clka; // @[util.scala 130:17]
  assign cluster_24_dina = io_dina; // @[util.scala 134:17]
  assign cluster_24_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_24_wea = io_wea & 18'h18 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_24_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_24_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_24_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_24_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_24_web = 1'h0; // @[util.scala 137:26]
  assign cluster_25_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_25_clka = io_clka; // @[util.scala 130:17]
  assign cluster_25_dina = io_dina; // @[util.scala 134:17]
  assign cluster_25_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_25_wea = io_wea & 18'h19 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_25_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_25_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_25_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_25_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_25_web = 1'h0; // @[util.scala 137:26]
  assign cluster_26_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_26_clka = io_clka; // @[util.scala 130:17]
  assign cluster_26_dina = io_dina; // @[util.scala 134:17]
  assign cluster_26_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_26_wea = io_wea & 18'h1a == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_26_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_26_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_26_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_26_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_26_web = 1'h0; // @[util.scala 137:26]
  assign cluster_27_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_27_clka = io_clka; // @[util.scala 130:17]
  assign cluster_27_dina = io_dina; // @[util.scala 134:17]
  assign cluster_27_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_27_wea = io_wea & 18'h1b == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_27_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_27_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_27_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_27_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_27_web = 1'h0; // @[util.scala 137:26]
  assign cluster_28_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_28_clka = io_clka; // @[util.scala 130:17]
  assign cluster_28_dina = io_dina; // @[util.scala 134:17]
  assign cluster_28_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_28_wea = io_wea & 18'h1c == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_28_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_28_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_28_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_28_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_28_web = 1'h0; // @[util.scala 137:26]
  assign cluster_29_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_29_clka = io_clka; // @[util.scala 130:17]
  assign cluster_29_dina = io_dina; // @[util.scala 134:17]
  assign cluster_29_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_29_wea = io_wea & 18'h1d == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_29_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_29_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_29_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_29_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_29_web = 1'h0; // @[util.scala 137:26]
  assign cluster_30_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_30_clka = io_clka; // @[util.scala 130:17]
  assign cluster_30_dina = io_dina; // @[util.scala 134:17]
  assign cluster_30_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_30_wea = io_wea & 18'h1e == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_30_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_30_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_30_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_30_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_30_web = 1'h0; // @[util.scala 137:26]
  assign cluster_31_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_31_clka = io_clka; // @[util.scala 130:17]
  assign cluster_31_dina = io_dina; // @[util.scala 134:17]
  assign cluster_31_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_31_wea = io_wea & 18'h1f == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_31_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_31_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_31_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_31_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_31_web = 1'h0; // @[util.scala 137:26]
  assign cluster_32_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_32_clka = io_clka; // @[util.scala 130:17]
  assign cluster_32_dina = io_dina; // @[util.scala 134:17]
  assign cluster_32_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_32_wea = io_wea & 18'h20 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_32_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_32_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_32_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_32_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_32_web = 1'h0; // @[util.scala 137:26]
  assign cluster_33_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_33_clka = io_clka; // @[util.scala 130:17]
  assign cluster_33_dina = io_dina; // @[util.scala 134:17]
  assign cluster_33_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_33_wea = io_wea & 18'h21 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_33_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_33_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_33_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_33_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_33_web = 1'h0; // @[util.scala 137:26]
  assign cluster_34_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_34_clka = io_clka; // @[util.scala 130:17]
  assign cluster_34_dina = io_dina; // @[util.scala 134:17]
  assign cluster_34_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_34_wea = io_wea & 18'h22 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_34_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_34_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_34_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_34_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_34_web = 1'h0; // @[util.scala 137:26]
  assign cluster_35_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_35_clka = io_clka; // @[util.scala 130:17]
  assign cluster_35_dina = io_dina; // @[util.scala 134:17]
  assign cluster_35_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_35_wea = io_wea & 18'h23 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_35_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_35_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_35_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_35_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_35_web = 1'h0; // @[util.scala 137:26]
  assign cluster_36_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_36_clka = io_clka; // @[util.scala 130:17]
  assign cluster_36_dina = io_dina; // @[util.scala 134:17]
  assign cluster_36_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_36_wea = io_wea & 18'h24 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_36_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_36_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_36_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_36_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_36_web = 1'h0; // @[util.scala 137:26]
  assign cluster_37_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_37_clka = io_clka; // @[util.scala 130:17]
  assign cluster_37_dina = io_dina; // @[util.scala 134:17]
  assign cluster_37_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_37_wea = io_wea & 18'h25 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_37_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_37_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_37_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_37_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_37_web = 1'h0; // @[util.scala 137:26]
  assign cluster_38_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_38_clka = io_clka; // @[util.scala 130:17]
  assign cluster_38_dina = io_dina; // @[util.scala 134:17]
  assign cluster_38_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_38_wea = io_wea & 18'h26 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_38_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_38_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_38_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_38_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_38_web = 1'h0; // @[util.scala 137:26]
  assign cluster_39_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_39_clka = io_clka; // @[util.scala 130:17]
  assign cluster_39_dina = io_dina; // @[util.scala 134:17]
  assign cluster_39_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_39_wea = io_wea & 18'h27 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_39_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_39_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_39_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_39_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_39_web = 1'h0; // @[util.scala 137:26]
  assign cluster_40_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_40_clka = io_clka; // @[util.scala 130:17]
  assign cluster_40_dina = io_dina; // @[util.scala 134:17]
  assign cluster_40_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_40_wea = io_wea & 18'h28 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_40_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_40_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_40_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_40_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_40_web = 1'h0; // @[util.scala 137:26]
  assign cluster_41_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_41_clka = io_clka; // @[util.scala 130:17]
  assign cluster_41_dina = io_dina; // @[util.scala 134:17]
  assign cluster_41_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_41_wea = io_wea & 18'h29 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_41_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_41_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_41_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_41_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_41_web = 1'h0; // @[util.scala 137:26]
  assign cluster_42_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_42_clka = io_clka; // @[util.scala 130:17]
  assign cluster_42_dina = io_dina; // @[util.scala 134:17]
  assign cluster_42_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_42_wea = io_wea & 18'h2a == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_42_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_42_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_42_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_42_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_42_web = 1'h0; // @[util.scala 137:26]
  assign cluster_43_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_43_clka = io_clka; // @[util.scala 130:17]
  assign cluster_43_dina = io_dina; // @[util.scala 134:17]
  assign cluster_43_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_43_wea = io_wea & 18'h2b == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_43_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_43_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_43_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_43_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_43_web = 1'h0; // @[util.scala 137:26]
  assign cluster_44_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_44_clka = io_clka; // @[util.scala 130:17]
  assign cluster_44_dina = io_dina; // @[util.scala 134:17]
  assign cluster_44_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_44_wea = io_wea & 18'h2c == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_44_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_44_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_44_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_44_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_44_web = 1'h0; // @[util.scala 137:26]
  assign cluster_45_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_45_clka = io_clka; // @[util.scala 130:17]
  assign cluster_45_dina = io_dina; // @[util.scala 134:17]
  assign cluster_45_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_45_wea = io_wea & 18'h2d == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_45_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_45_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_45_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_45_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_45_web = 1'h0; // @[util.scala 137:26]
  assign cluster_46_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_46_clka = io_clka; // @[util.scala 130:17]
  assign cluster_46_dina = io_dina; // @[util.scala 134:17]
  assign cluster_46_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_46_wea = io_wea & 18'h2e == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_46_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_46_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_46_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_46_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_46_web = 1'h0; // @[util.scala 137:26]
  assign cluster_47_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_47_clka = io_clka; // @[util.scala 130:17]
  assign cluster_47_dina = io_dina; // @[util.scala 134:17]
  assign cluster_47_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_47_wea = io_wea & 18'h2f == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_47_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_47_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_47_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_47_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_47_web = 1'h0; // @[util.scala 137:26]
  assign cluster_48_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_48_clka = io_clka; // @[util.scala 130:17]
  assign cluster_48_dina = io_dina; // @[util.scala 134:17]
  assign cluster_48_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_48_wea = io_wea & 18'h30 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_48_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_48_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_48_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_48_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_48_web = 1'h0; // @[util.scala 137:26]
  assign cluster_49_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_49_clka = io_clka; // @[util.scala 130:17]
  assign cluster_49_dina = io_dina; // @[util.scala 134:17]
  assign cluster_49_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_49_wea = io_wea & 18'h31 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_49_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_49_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_49_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_49_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_49_web = 1'h0; // @[util.scala 137:26]
  assign cluster_50_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_50_clka = io_clka; // @[util.scala 130:17]
  assign cluster_50_dina = io_dina; // @[util.scala 134:17]
  assign cluster_50_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_50_wea = io_wea & 18'h32 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_50_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_50_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_50_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_50_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_50_web = 1'h0; // @[util.scala 137:26]
  assign cluster_51_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_51_clka = io_clka; // @[util.scala 130:17]
  assign cluster_51_dina = io_dina; // @[util.scala 134:17]
  assign cluster_51_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_51_wea = io_wea & 18'h33 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_51_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_51_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_51_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_51_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_51_web = 1'h0; // @[util.scala 137:26]
  assign cluster_52_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_52_clka = io_clka; // @[util.scala 130:17]
  assign cluster_52_dina = io_dina; // @[util.scala 134:17]
  assign cluster_52_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_52_wea = io_wea & 18'h34 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_52_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_52_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_52_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_52_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_52_web = 1'h0; // @[util.scala 137:26]
  assign cluster_53_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_53_clka = io_clka; // @[util.scala 130:17]
  assign cluster_53_dina = io_dina; // @[util.scala 134:17]
  assign cluster_53_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_53_wea = io_wea & 18'h35 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_53_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_53_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_53_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_53_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_53_web = 1'h0; // @[util.scala 137:26]
  assign cluster_54_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_54_clka = io_clka; // @[util.scala 130:17]
  assign cluster_54_dina = io_dina; // @[util.scala 134:17]
  assign cluster_54_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_54_wea = io_wea & 18'h36 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_54_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_54_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_54_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_54_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_54_web = 1'h0; // @[util.scala 137:26]
  assign cluster_55_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_55_clka = io_clka; // @[util.scala 130:17]
  assign cluster_55_dina = io_dina; // @[util.scala 134:17]
  assign cluster_55_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_55_wea = io_wea & 18'h37 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_55_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_55_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_55_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_55_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_55_web = 1'h0; // @[util.scala 137:26]
  assign cluster_56_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_56_clka = io_clka; // @[util.scala 130:17]
  assign cluster_56_dina = io_dina; // @[util.scala 134:17]
  assign cluster_56_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_56_wea = io_wea & 18'h38 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_56_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_56_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_56_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_56_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_56_web = 1'h0; // @[util.scala 137:26]
  assign cluster_57_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_57_clka = io_clka; // @[util.scala 130:17]
  assign cluster_57_dina = io_dina; // @[util.scala 134:17]
  assign cluster_57_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_57_wea = io_wea & 18'h39 == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_57_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_57_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_57_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_57_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_57_web = 1'h0; // @[util.scala 137:26]
  assign cluster_58_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_58_clka = io_clka; // @[util.scala 130:17]
  assign cluster_58_dina = io_dina; // @[util.scala 134:17]
  assign cluster_58_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_58_wea = io_wea & 18'h3a == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_58_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_58_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_58_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_58_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_58_web = 1'h0; // @[util.scala 137:26]
  assign cluster_59_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_59_clka = io_clka; // @[util.scala 130:17]
  assign cluster_59_dina = io_dina; // @[util.scala 134:17]
  assign cluster_59_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_59_wea = io_wea & 18'h3b == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_59_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_59_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_59_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_59_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_59_web = 1'h0; // @[util.scala 137:26]
  assign cluster_60_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_60_clka = io_clka; // @[util.scala 130:17]
  assign cluster_60_dina = io_dina; // @[util.scala 134:17]
  assign cluster_60_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_60_wea = io_wea & 18'h3c == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_60_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_60_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_60_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_60_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_60_web = 1'h0; // @[util.scala 137:26]
  assign cluster_61_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_61_clka = io_clka; // @[util.scala 130:17]
  assign cluster_61_dina = io_dina; // @[util.scala 134:17]
  assign cluster_61_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_61_wea = io_wea & 18'h3d == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_61_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_61_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_61_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_61_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_61_web = 1'h0; // @[util.scala 137:26]
  assign cluster_62_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_62_clka = io_clka; // @[util.scala 130:17]
  assign cluster_62_dina = io_dina; // @[util.scala 134:17]
  assign cluster_62_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_62_wea = io_wea & 18'h3e == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_62_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_62_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_62_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_62_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_62_web = 1'h0; // @[util.scala 137:26]
  assign cluster_63_addra = io_addra[11:0]; // @[util.scala 136:29]
  assign cluster_63_clka = io_clka; // @[util.scala 130:17]
  assign cluster_63_dina = io_dina; // @[util.scala 134:17]
  assign cluster_63_ena = 1'h1; // @[util.scala 132:16]
  assign cluster_63_wea = io_wea & 18'h3f == _cluster_0_io_wea_T; // @[util.scala 138:26]
  assign cluster_63_addrb = io_addrb[11:0]; // @[util.scala 135:29]
  assign cluster_63_clkb = io_clkb; // @[util.scala 129:17]
  assign cluster_63_dinb = 48'h0; // @[util.scala 133:17]
  assign cluster_63_enb = 1'h1; // @[util.scala 131:16]
  assign cluster_63_web = 1'h0; // @[util.scala 137:26]
endmodule
module pipeline_97(
  input         clock,
  input         reset,
  input         io_dout_ready,
  output        io_dout_valid,
  output [15:0] io_dout_bits_addr,
  output [11:0] io_dout_bits_block_index,
  output        io_din_ready,
  input         io_din_valid,
  input  [15:0] io_din_bits_addr,
  input  [11:0] io_din_bits_block_index
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] data_addr; // @[util.scala 238:21]
  reg [11:0] data_block_index; // @[util.scala 238:21]
  reg  valid; // @[util.scala 239:22]
  reg  ready; // @[util.scala 240:22]
  reg [15:0] data2_addr; // @[util.scala 241:22]
  reg [11:0] data2_block_index; // @[util.scala 241:22]
  reg  valid2; // @[util.scala 242:23]
  wire  _GEN_2 = ready & io_din_valid; // @[util.scala 247:22 util.scala 249:13 util.scala 252:13]
  assign io_dout_valid = valid; // @[util.scala 268:17]
  assign io_dout_bits_addr = data_addr; // @[util.scala 269:16]
  assign io_dout_bits_block_index = data_block_index; // @[util.scala 269:16]
  assign io_din_ready = ready; // @[util.scala 267:16]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 238:21]
      data_addr <= 16'h0; // @[util.scala 238:21]
    end else if (io_dout_ready) begin // @[util.scala 243:22]
      if (valid2) begin // @[util.scala 244:17]
        data_addr <= data2_addr; // @[util.scala 245:12]
      end else if (ready) begin // @[util.scala 247:22]
        data_addr <= io_din_bits_addr; // @[util.scala 248:12]
      end else begin
        data_addr <= 16'h0; // @[util.scala 251:12]
      end
    end
    if (reset) begin // @[util.scala 238:21]
      data_block_index <= 12'h0; // @[util.scala 238:21]
    end else if (io_dout_ready) begin // @[util.scala 243:22]
      if (valid2) begin // @[util.scala 244:17]
        data_block_index <= data2_block_index; // @[util.scala 245:12]
      end else if (ready) begin // @[util.scala 247:22]
        data_block_index <= io_din_bits_block_index; // @[util.scala 248:12]
      end else begin
        data_block_index <= 12'h0; // @[util.scala 251:12]
      end
    end
    if (reset) begin // @[util.scala 239:22]
      valid <= 1'h0; // @[util.scala 239:22]
    end else if (io_dout_ready) begin // @[util.scala 243:22]
      if (valid2) begin // @[util.scala 244:17]
        valid <= valid2; // @[util.scala 246:13]
      end else begin
        valid <= _GEN_2;
      end
    end
    if (reset) begin // @[util.scala 240:22]
      ready <= 1'h0; // @[util.scala 240:22]
    end else begin
      ready <= io_dout_ready; // @[util.scala 255:9]
    end
    if (reset) begin // @[util.scala 241:22]
      data2_addr <= 16'h0; // @[util.scala 241:22]
    end else if (~io_dout_ready & ready) begin // @[util.scala 258:33]
      data2_addr <= io_din_bits_addr; // @[util.scala 259:11]
    end else if (io_dout_ready) begin // @[util.scala 261:28]
      data2_addr <= 16'h0; // @[util.scala 263:11]
    end
    if (reset) begin // @[util.scala 241:22]
      data2_block_index <= 12'h0; // @[util.scala 241:22]
    end else if (~io_dout_ready & ready) begin // @[util.scala 258:33]
      data2_block_index <= io_din_bits_block_index; // @[util.scala 259:11]
    end else if (io_dout_ready) begin // @[util.scala 261:28]
      data2_block_index <= 12'h0; // @[util.scala 263:11]
    end
    if (reset) begin // @[util.scala 242:23]
      valid2 <= 1'h0; // @[util.scala 242:23]
    end else if (~io_dout_ready & ready) begin // @[util.scala 258:33]
      valid2 <= io_din_valid; // @[util.scala 260:12]
    end else if (io_dout_ready) begin // @[util.scala 261:28]
      valid2 <= 1'h0; // @[util.scala 264:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_addr = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  data_block_index = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ready = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  data2_addr = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  data2_block_index = _RAND_5[11:0];
  _RAND_6 = {1{`RANDOM}};
  valid2 = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WB_engine(
  input          clock,
  input          reset,
  input          io_ddr_aw_ready,
  output         io_ddr_aw_valid,
  output [63:0]  io_ddr_aw_bits_awaddr,
  output [6:0]   io_ddr_aw_bits_awid,
  input          io_ddr_w_ready,
  output         io_ddr_w_valid,
  output [511:0] io_ddr_w_bits_wdata,
  output [63:0]  io_ddr_w_bits_wstrb,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [31:0]  io_xbar_in_bits_tdata,
  input  [63:0]  io_level_base_addr,
  input  [31:0]  io_level,
  output         io_end,
  input          io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [17:0] buffer_io_addra; // @[BFS.scala 23:22]
  wire  buffer_io_clka; // @[BFS.scala 23:22]
  wire [47:0] buffer_io_dina; // @[BFS.scala 23:22]
  wire  buffer_io_wea; // @[BFS.scala 23:22]
  wire [17:0] buffer_io_addrb; // @[BFS.scala 23:22]
  wire  buffer_io_clkb; // @[BFS.scala 23:22]
  wire [47:0] buffer_io_doutb; // @[BFS.scala 23:22]
  wire [11:0] region_counter__addra; // @[BFS.scala 24:30]
  wire  region_counter__clka; // @[BFS.scala 24:30]
  wire [8:0] region_counter__dina; // @[BFS.scala 24:30]
  wire  region_counter__ena; // @[BFS.scala 24:30]
  wire  region_counter__wea; // @[BFS.scala 24:30]
  wire [11:0] region_counter__addrb; // @[BFS.scala 24:30]
  wire  region_counter__clkb; // @[BFS.scala 24:30]
  wire [8:0] region_counter__doutb; // @[BFS.scala 24:30]
  wire  region_counter__enb; // @[BFS.scala 24:30]
  wire  region_counter_doutb_forward_clock; // @[BFS.scala 47:44]
  wire  region_counter_doutb_forward_reset; // @[BFS.scala 47:44]
  wire  region_counter_doutb_forward_io_dout_ready; // @[BFS.scala 47:44]
  wire  region_counter_doutb_forward_io_dout_valid; // @[BFS.scala 47:44]
  wire [8:0] region_counter_doutb_forward_io_dout_bits; // @[BFS.scala 47:44]
  wire  region_counter_doutb_forward_io_din_valid; // @[BFS.scala 47:44]
  wire [8:0] region_counter_doutb_forward_io_din_bits; // @[BFS.scala 47:44]
  wire  pipeline_1_clock; // @[BFS.scala 49:26]
  wire  pipeline_1_reset; // @[BFS.scala 49:26]
  wire  pipeline_1_io_dout_ready; // @[BFS.scala 49:26]
  wire  pipeline_1_io_dout_valid; // @[BFS.scala 49:26]
  wire [15:0] pipeline_1_io_dout_bits_addr; // @[BFS.scala 49:26]
  wire [11:0] pipeline_1_io_dout_bits_block_index; // @[BFS.scala 49:26]
  wire  pipeline_1_io_din_ready; // @[BFS.scala 49:26]
  wire  pipeline_1_io_din_valid; // @[BFS.scala 49:26]
  wire [15:0] pipeline_1_io_din_bits_addr; // @[BFS.scala 49:26]
  wire [11:0] pipeline_1_io_din_bits_block_index; // @[BFS.scala 49:26]
  wire  aw_buffer_full; // @[BFS.scala 82:25]
  wire [63:0] aw_buffer_din; // @[BFS.scala 82:25]
  wire  aw_buffer_wr_en; // @[BFS.scala 82:25]
  wire  aw_buffer_empty; // @[BFS.scala 82:25]
  wire [63:0] aw_buffer_dout; // @[BFS.scala 82:25]
  wire  aw_buffer_rd_en; // @[BFS.scala 82:25]
  wire [5:0] aw_buffer_data_count; // @[BFS.scala 82:25]
  wire  aw_buffer_clk; // @[BFS.scala 82:25]
  wire  aw_buffer_srst; // @[BFS.scala 82:25]
  wire  aw_buffer_valid; // @[BFS.scala 82:25]
  wire  w_buffer_full; // @[BFS.scala 83:24]
  wire [63:0] w_buffer_din; // @[BFS.scala 83:24]
  wire  w_buffer_wr_en; // @[BFS.scala 83:24]
  wire  w_buffer_empty; // @[BFS.scala 83:24]
  wire [63:0] w_buffer_dout; // @[BFS.scala 83:24]
  wire  w_buffer_rd_en; // @[BFS.scala 83:24]
  wire [5:0] w_buffer_data_count; // @[BFS.scala 83:24]
  wire  w_buffer_clk; // @[BFS.scala 83:24]
  wire  w_buffer_srst; // @[BFS.scala 83:24]
  wire  w_buffer_valid; // @[BFS.scala 83:24]
  wire [33:0] _GEN_16 = {io_xbar_in_bits_tdata, 2'h0}; // @[BFS.scala 37:23]
  wire [34:0] _dramaddr_T = {{1'd0}, _GEN_16}; // @[BFS.scala 37:23]
  wire [63:0] dramaddr = {{29'd0}, _dramaddr_T}; // @[BFS.scala 37:39 BFS.scala 37:39]
  wire [11:0] block_index = dramaddr[25:14]; // @[BFS.scala 38:29]
  wire  _pipeline_1_io_din_valid_T = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 53:47]
  wire  _buffer_io_wea_T = pipeline_1_io_dout_valid & pipeline_1_io_dout_ready; // @[BFS.scala 59:45]
  wire [8:0] region_counter_doutb = region_counter_doutb_forward_io_dout_valid ?
    region_counter_doutb_forward_io_dout_bits : region_counter__doutb; // @[BFS.scala 71:30]
  wire [5:0] buffer_io_addra_lo = region_counter_doutb[5:0]; // @[BFS.scala 27:35 BFS.scala 27:35]
  wire  _region_counter_dina_0_T = region_counter_doutb == 9'h3f; // @[BFS.scala 31:17]
  wire [8:0] _region_counter_dina_0_T_2 = region_counter_doutb + 9'h1; // @[BFS.scala 31:40]
  wire [8:0] region_counter_dina_0 = region_counter_doutb == 9'h3f ? 9'h0 : _region_counter_dina_0_T_2; // @[BFS.scala 31:8]
  wire  _region_counter_doutb_forward_io_din_valid_T_1 = pipeline_1_io_dout_bits_block_index == block_index; // @[BFS.scala 69:28]
  wire  _region_counter_doutb_forward_io_din_valid_T_2 = _pipeline_1_io_din_valid_T &
    _region_counter_doutb_forward_io_din_valid_T_1; // @[BFS.scala 68:85]
  reg [1:0] wb_sm; // @[BFS.scala 80:22]
  reg [7:0] count; // @[BFS.scala 81:22]
  reg [11:0] wb_block_index; // @[BFS.scala 84:31]
  wire  _flush_start_T = wb_sm == 2'h0; // @[BFS.scala 85:28]
  wire  flush_start = wb_sm == 2'h0 & io_flush; // @[BFS.scala 85:42]
  reg [7:0] size_b; // @[BFS.scala 86:23]
  reg [63:0] level_base_addr_reg; // @[BFS.scala 87:36]
  wire  wb_start = pipeline_1_io_dout_valid & _region_counter_dina_0_T & _flush_start_T; // @[BFS.scala 88:77]
  wire  _T = wb_sm == 2'h3; // @[BFS.scala 95:20]
  wire [8:0] _GEN_0 = wb_sm == 2'h3 ? region_counter_doutb : {{1'd0}, size_b}; // @[BFS.scala 95:38 BFS.scala 96:12 BFS.scala 86:23]
  wire [8:0] _GEN_1 = wb_start ? 9'h40 : _GEN_0; // @[BFS.scala 93:17 BFS.scala 94:12]
  wire  _T_1 = wb_sm == 2'h2; // @[BFS.scala 103:20]
  wire  _T_2 = wb_block_index != 12'hfff; // @[BFS.scala 103:55]
  wire [11:0] _wb_block_index_T_1 = wb_block_index + 12'h1; // @[BFS.scala 104:38]
  wire  _T_6 = wb_sm == 2'h1; // @[BFS.scala 118:20]
  wire  _T_7 = ~aw_buffer_full; // @[BFS.scala 118:57]
  wire  _T_9 = ~w_buffer_full; // @[BFS.scala 118:89]
  wire  _T_10 = wb_sm == 2'h1 & ~aw_buffer_full & ~w_buffer_full; // @[BFS.scala 118:69]
  wire [1:0] _GEN_6 = io_flush ? 2'h2 : 2'h0; // @[BFS.scala 120:21 BFS.scala 121:15 BFS.scala 123:15]
  wire [1:0] _GEN_7 = count == size_b ? _GEN_6 : 2'h1; // @[BFS.scala 119:27 BFS.scala 126:13]
  wire [1:0] _GEN_8 = _T_2 ? 2'h3 : 2'h0; // @[BFS.scala 129:46 BFS.scala 130:13 BFS.scala 132:13]
  wire [1:0] _GEN_9 = _T_1 ? _GEN_8 : wb_sm; // @[BFS.scala 128:38 BFS.scala 80:22]
  wire [1:0] _GEN_10 = wb_sm == 2'h1 & ~aw_buffer_full & ~w_buffer_full ? _GEN_7 : _GEN_9; // @[BFS.scala 118:102]
  wire [7:0] _count_T_1 = count + 8'h1; // @[BFS.scala 139:20]
  wire [17:0] _buffer_io_addrb_T = {block_index,6'h0}; // @[Cat.scala 30:58]
  wire [5:0] buffer_io_addrb_lo_2 = count[5:0]; // @[BFS.scala 27:35 BFS.scala 27:35]
  wire [17:0] _buffer_io_addrb_T_4 = {wb_block_index,buffer_io_addrb_lo_2}; // @[Cat.scala 30:58]
  wire [17:0] _buffer_io_addrb_T_5 = wb_start ? _buffer_io_addrb_T : 18'h0; // @[Mux.scala 27:72]
  wire [17:0] _buffer_io_addrb_T_6 = _T ? _buffer_io_addrb_T : 18'h0; // @[Mux.scala 27:72]
  wire [17:0] _buffer_io_addrb_T_7 = _T_6 ? _buffer_io_addrb_T_4 : 18'h0; // @[Mux.scala 27:72]
  wire [17:0] _buffer_io_addrb_T_8 = _buffer_io_addrb_T_5 | _buffer_io_addrb_T_6; // @[Mux.scala 27:72]
  wire [11:0] _region_counter_io_addrb_T_4 = _T_6 ? pipeline_1_io_dout_bits_block_index : block_index; // @[Mux.scala 98:16]
  wire [11:0] _region_counter_io_addrb_T_5 = flush_start ? 12'h0 : _region_counter_io_addrb_T_4; // @[Mux.scala 98:16]
  wire [13:0] aw_buffer_io_din_lo = buffer_io_doutb[45:32]; // @[BFS.scala 164:80]
  wire [25:0] _aw_buffer_io_din_T = {wb_block_index,aw_buffer_io_din_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_17 = {{38'd0}, _aw_buffer_io_din_T}; // @[BFS.scala 164:43]
  wire [57:0] alignment_addr = aw_buffer_dout[63:6]; // @[BFS.scala 165:41]
  wire [5:0] io_ddr_aw_bits_awid_lo = aw_buffer_data_count; // @[BFS.scala 168:72 BFS.scala 168:72]
  wire [5:0] alignment_offset = w_buffer_dout[37:32]; // @[BFS.scala 179:42]
  wire [9:0] _io_ddr_w_bits_wdata_T_1 = 4'h8 * alignment_offset; // @[BFS.scala 180:80]
  wire [511:0] _io_ddr_w_bits_wdata_WIRE = {{480'd0}, w_buffer_dout[31:0]}; // @[BFS.scala 180:58 BFS.scala 180:58]
  wire [1534:0] _GEN_18 = {{1023'd0}, _io_ddr_w_bits_wdata_WIRE}; // @[BFS.scala 180:72]
  wire [1534:0] _io_ddr_w_bits_wdata_T_2 = _GEN_18 << _io_ddr_w_bits_wdata_T_1; // @[BFS.scala 180:72]
  wire [126:0] _io_ddr_w_bits_wstrb_T = 127'hf << alignment_offset; // @[BFS.scala 183:38]
  URAM_cluster buffer ( // @[BFS.scala 23:22]
    .io_addra(buffer_io_addra),
    .io_clka(buffer_io_clka),
    .io_dina(buffer_io_dina),
    .io_wea(buffer_io_wea),
    .io_addrb(buffer_io_addrb),
    .io_clkb(buffer_io_clkb),
    .io_doutb(buffer_io_doutb)
  );
  region_counter region_counter_ ( // @[BFS.scala 24:30]
    .addra(region_counter__addra),
    .clka(region_counter__clka),
    .dina(region_counter__dina),
    .ena(region_counter__ena),
    .wea(region_counter__wea),
    .addrb(region_counter__addrb),
    .clkb(region_counter__clkb),
    .doutb(region_counter__doutb),
    .enb(region_counter__enb)
  );
  pipeline_34 region_counter_doutb_forward ( // @[BFS.scala 47:44]
    .clock(region_counter_doutb_forward_clock),
    .reset(region_counter_doutb_forward_reset),
    .io_dout_ready(region_counter_doutb_forward_io_dout_ready),
    .io_dout_valid(region_counter_doutb_forward_io_dout_valid),
    .io_dout_bits(region_counter_doutb_forward_io_dout_bits),
    .io_din_valid(region_counter_doutb_forward_io_din_valid),
    .io_din_bits(region_counter_doutb_forward_io_din_bits)
  );
  pipeline_97 pipeline_1 ( // @[BFS.scala 49:26]
    .clock(pipeline_1_clock),
    .reset(pipeline_1_reset),
    .io_dout_ready(pipeline_1_io_dout_ready),
    .io_dout_valid(pipeline_1_io_dout_valid),
    .io_dout_bits_addr(pipeline_1_io_dout_bits_addr),
    .io_dout_bits_block_index(pipeline_1_io_dout_bits_block_index),
    .io_din_ready(pipeline_1_io_din_ready),
    .io_din_valid(pipeline_1_io_din_valid),
    .io_din_bits_addr(pipeline_1_io_din_bits_addr),
    .io_din_bits_block_index(pipeline_1_io_din_bits_block_index)
  );
  addr_fifo aw_buffer ( // @[BFS.scala 82:25]
    .full(aw_buffer_full),
    .din(aw_buffer_din),
    .wr_en(aw_buffer_wr_en),
    .empty(aw_buffer_empty),
    .dout(aw_buffer_dout),
    .rd_en(aw_buffer_rd_en),
    .data_count(aw_buffer_data_count),
    .clk(aw_buffer_clk),
    .srst(aw_buffer_srst),
    .valid(aw_buffer_valid)
  );
  level_fifo w_buffer ( // @[BFS.scala 83:24]
    .full(w_buffer_full),
    .din(w_buffer_din),
    .wr_en(w_buffer_wr_en),
    .empty(w_buffer_empty),
    .dout(w_buffer_dout),
    .rd_en(w_buffer_rd_en),
    .data_count(w_buffer_data_count),
    .clk(w_buffer_clk),
    .srst(w_buffer_srst),
    .valid(w_buffer_valid)
  );
  assign io_ddr_aw_valid = aw_buffer_valid; // @[BFS.scala 172:19]
  assign io_ddr_aw_bits_awaddr = {alignment_addr,6'h0}; // @[Cat.scala 30:58]
  assign io_ddr_aw_bits_awid = {1'h1,io_ddr_aw_bits_awid_lo}; // @[Cat.scala 30:58]
  assign io_ddr_w_valid = w_buffer_valid; // @[BFS.scala 182:18]
  assign io_ddr_w_bits_wdata = _io_ddr_w_bits_wdata_T_2[511:0]; // @[BFS.scala 180:23]
  assign io_ddr_w_bits_wstrb = _io_ddr_w_bits_wstrb_T[63:0]; // @[BFS.scala 183:23]
  assign io_xbar_in_ready = pipeline_1_io_din_ready; // @[BFS.scala 56:20]
  assign io_end = _T_1 & wb_block_index == 12'hfff; // @[BFS.scala 188:36]
  assign buffer_io_addra = {pipeline_1_io_dout_bits_block_index,buffer_io_addra_lo}; // @[Cat.scala 30:58]
  assign buffer_io_clka = clock; // @[BFS.scala 62:33]
  assign buffer_io_dina = {pipeline_1_io_dout_bits_addr,io_level}; // @[Cat.scala 30:58]
  assign buffer_io_wea = pipeline_1_io_dout_valid & pipeline_1_io_dout_ready; // @[BFS.scala 59:45]
  assign buffer_io_addrb = _buffer_io_addrb_T_8 | _buffer_io_addrb_T_7; // @[Mux.scala 27:72]
  assign buffer_io_clkb = clock; // @[BFS.scala 150:33]
  assign region_counter__addra = _T_6 ? wb_block_index : pipeline_1_io_dout_bits_block_index; // @[BFS.scala 152:33]
  assign region_counter__clka = clock; // @[BFS.scala 41:41]
  assign region_counter__dina = _T_6 ? 9'h0 : region_counter_dina_0; // @[BFS.scala 154:32]
  assign region_counter__ena = 1'h1; // @[BFS.scala 42:25]
  assign region_counter__wea = _T_6 | _buffer_io_wea_T; // @[BFS.scala 153:31]
  assign region_counter__addrb = _T_1 ? _wb_block_index_T_1 : _region_counter_io_addrb_T_5; // @[Mux.scala 98:16]
  assign region_counter__clkb = clock; // @[BFS.scala 40:41]
  assign region_counter__enb = 1'h1; // @[BFS.scala 43:25]
  assign region_counter_doutb_forward_clock = clock;
  assign region_counter_doutb_forward_reset = reset;
  assign region_counter_doutb_forward_io_dout_ready = wb_sm == 2'h0; // @[BFS.scala 90:55]
  assign region_counter_doutb_forward_io_din_valid = _region_counter_doutb_forward_io_din_valid_T_2 & _buffer_io_wea_T; // @[BFS.scala 69:55]
  assign region_counter_doutb_forward_io_din_bits = region_counter_doutb == 9'h3f ? 9'h0 : _region_counter_dina_0_T_2; // @[BFS.scala 31:8]
  assign pipeline_1_clock = clock;
  assign pipeline_1_reset = reset;
  assign pipeline_1_io_dout_ready = wb_sm == 2'h0; // @[BFS.scala 89:37]
  assign pipeline_1_io_din_valid = io_xbar_in_valid & io_xbar_in_ready; // @[BFS.scala 53:47]
  assign pipeline_1_io_din_bits_addr = {{2'd0}, dramaddr[13:0]}; // @[BFS.scala 54:58 BFS.scala 54:58]
  assign pipeline_1_io_din_bits_block_index = dramaddr[25:14]; // @[BFS.scala 38:29]
  assign aw_buffer_din = level_base_addr_reg + _GEN_17; // @[BFS.scala 164:43]
  assign aw_buffer_wr_en = _T_6 & _T_9; // @[BFS.scala 163:47]
  assign aw_buffer_rd_en = io_ddr_aw_ready; // @[BFS.scala 173:22]
  assign aw_buffer_clk = clock; // @[BFS.scala 161:35]
  assign aw_buffer_srst = reset; // @[BFS.scala 162:36]
  assign w_buffer_din = {{26'd0}, buffer_io_doutb[37:0]}; // @[BFS.scala 178:37]
  assign w_buffer_wr_en = _T_6 & _T_7; // @[BFS.scala 177:46]
  assign w_buffer_rd_en = io_ddr_w_ready; // @[BFS.scala 184:21]
  assign w_buffer_clk = clock; // @[BFS.scala 175:34]
  assign w_buffer_srst = reset; // @[BFS.scala 176:35]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 80:22]
      wb_sm <= 2'h0; // @[BFS.scala 80:22]
    end else if (flush_start) begin // @[BFS.scala 108:20]
      wb_sm <= 2'h3; // @[BFS.scala 109:11]
    end else if (_T) begin // @[BFS.scala 110:38]
      if (region_counter_doutb == 9'h0) begin // @[BFS.scala 111:39]
        wb_sm <= 2'h2; // @[BFS.scala 112:13]
      end else begin
        wb_sm <= 2'h1; // @[BFS.scala 114:13]
      end
    end else if (wb_start) begin // @[BFS.scala 116:23]
      wb_sm <= 2'h1; // @[BFS.scala 117:11]
    end else begin
      wb_sm <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 81:22]
      count <= 8'h0; // @[BFS.scala 81:22]
    end else if (_flush_start_T | _T_1) begin // @[BFS.scala 136:53]
      count <= 8'h1; // @[BFS.scala 137:11]
    end else if (_T_10) begin // @[BFS.scala 138:101]
      count <= _count_T_1; // @[BFS.scala 139:11]
    end
    if (reset) begin // @[BFS.scala 84:31]
      wb_block_index <= 12'h0; // @[BFS.scala 84:31]
    end else if (wb_start) begin // @[BFS.scala 99:17]
      wb_block_index <= pipeline_1_io_dout_bits_block_index; // @[BFS.scala 100:20]
    end else if (flush_start) begin // @[BFS.scala 101:26]
      wb_block_index <= 12'h0; // @[BFS.scala 102:20]
    end else if (wb_sm == 2'h2 & wb_block_index != 12'hfff) begin // @[BFS.scala 103:76]
      wb_block_index <= _wb_block_index_T_1; // @[BFS.scala 104:20]
    end
    if (reset) begin // @[BFS.scala 86:23]
      size_b <= 8'h0; // @[BFS.scala 86:23]
    end else begin
      size_b <= _GEN_1[7:0];
    end
    if (reset) begin // @[BFS.scala 87:36]
      level_base_addr_reg <= 64'h0; // @[BFS.scala 87:36]
    end else begin
      level_base_addr_reg <= io_level_base_addr; // @[BFS.scala 91:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_sm = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  wb_block_index = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  size_b = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  level_base_addr_reg = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Apply(
  input          clock,
  input          reset,
  input          io_ddr_aw_ready,
  output         io_ddr_aw_valid,
  output [63:0]  io_ddr_aw_bits_awaddr,
  output [6:0]   io_ddr_aw_bits_awid,
  input          io_ddr_w_ready,
  output         io_ddr_w_valid,
  output [511:0] io_ddr_w_bits_wdata,
  output [63:0]  io_ddr_w_bits_wstrb,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input  [31:0]  io_level,
  input  [63:0]  io_level_base_addr,
  output         io_end,
  input          io_flush
);
  wire  vertex_update_buffer_full; // @[BFS.scala 208:36]
  wire [63:0] vertex_update_buffer_din; // @[BFS.scala 208:36]
  wire  vertex_update_buffer_wr_en; // @[BFS.scala 208:36]
  wire  vertex_update_buffer_empty; // @[BFS.scala 208:36]
  wire [63:0] vertex_update_buffer_dout; // @[BFS.scala 208:36]
  wire  vertex_update_buffer_rd_en; // @[BFS.scala 208:36]
  wire [5:0] vertex_update_buffer_data_count; // @[BFS.scala 208:36]
  wire  vertex_update_buffer_clk; // @[BFS.scala 208:36]
  wire  vertex_update_buffer_srst; // @[BFS.scala 208:36]
  wire  vertex_update_buffer_valid; // @[BFS.scala 208:36]
  wire  update_engine_clock; // @[BFS.scala 217:29]
  wire  update_engine_reset; // @[BFS.scala 217:29]
  wire  update_engine_io_ddr_aw_ready; // @[BFS.scala 217:29]
  wire  update_engine_io_ddr_aw_valid; // @[BFS.scala 217:29]
  wire [63:0] update_engine_io_ddr_aw_bits_awaddr; // @[BFS.scala 217:29]
  wire [6:0] update_engine_io_ddr_aw_bits_awid; // @[BFS.scala 217:29]
  wire  update_engine_io_ddr_w_ready; // @[BFS.scala 217:29]
  wire  update_engine_io_ddr_w_valid; // @[BFS.scala 217:29]
  wire [511:0] update_engine_io_ddr_w_bits_wdata; // @[BFS.scala 217:29]
  wire [63:0] update_engine_io_ddr_w_bits_wstrb; // @[BFS.scala 217:29]
  wire  update_engine_io_xbar_in_ready; // @[BFS.scala 217:29]
  wire  update_engine_io_xbar_in_valid; // @[BFS.scala 217:29]
  wire [31:0] update_engine_io_xbar_in_bits_tdata; // @[BFS.scala 217:29]
  wire [63:0] update_engine_io_level_base_addr; // @[BFS.scala 217:29]
  wire [31:0] update_engine_io_level; // @[BFS.scala 217:29]
  wire  update_engine_io_end; // @[BFS.scala 217:29]
  wire  update_engine_io_flush; // @[BFS.scala 217:29]
  wire  FIN = io_gather_in_bits_tdata[31] & io_gather_in_valid; // @[BFS.scala 209:41]
  wire  _update_engine_io_flush_T = vertex_update_buffer_data_count == 6'h0; // @[util.scala 211:19]
  update_fifo vertex_update_buffer ( // @[BFS.scala 208:36]
    .full(vertex_update_buffer_full),
    .din(vertex_update_buffer_din),
    .wr_en(vertex_update_buffer_wr_en),
    .empty(vertex_update_buffer_empty),
    .dout(vertex_update_buffer_dout),
    .rd_en(vertex_update_buffer_rd_en),
    .data_count(vertex_update_buffer_data_count),
    .clk(vertex_update_buffer_clk),
    .srst(vertex_update_buffer_srst),
    .valid(vertex_update_buffer_valid)
  );
  WB_engine update_engine ( // @[BFS.scala 217:29]
    .clock(update_engine_clock),
    .reset(update_engine_reset),
    .io_ddr_aw_ready(update_engine_io_ddr_aw_ready),
    .io_ddr_aw_valid(update_engine_io_ddr_aw_valid),
    .io_ddr_aw_bits_awaddr(update_engine_io_ddr_aw_bits_awaddr),
    .io_ddr_aw_bits_awid(update_engine_io_ddr_aw_bits_awid),
    .io_ddr_w_ready(update_engine_io_ddr_w_ready),
    .io_ddr_w_valid(update_engine_io_ddr_w_valid),
    .io_ddr_w_bits_wdata(update_engine_io_ddr_w_bits_wdata),
    .io_ddr_w_bits_wstrb(update_engine_io_ddr_w_bits_wstrb),
    .io_xbar_in_ready(update_engine_io_xbar_in_ready),
    .io_xbar_in_valid(update_engine_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(update_engine_io_xbar_in_bits_tdata),
    .io_level_base_addr(update_engine_io_level_base_addr),
    .io_level(update_engine_io_level),
    .io_end(update_engine_io_end),
    .io_flush(update_engine_io_flush)
  );
  assign io_ddr_aw_valid = update_engine_io_ddr_aw_valid; // @[BFS.scala 227:13]
  assign io_ddr_aw_bits_awaddr = update_engine_io_ddr_aw_bits_awaddr; // @[BFS.scala 227:13]
  assign io_ddr_aw_bits_awid = update_engine_io_ddr_aw_bits_awid; // @[BFS.scala 227:13]
  assign io_ddr_w_valid = update_engine_io_ddr_w_valid; // @[BFS.scala 228:12]
  assign io_ddr_w_bits_wdata = update_engine_io_ddr_w_bits_wdata; // @[BFS.scala 228:12]
  assign io_ddr_w_bits_wstrb = update_engine_io_ddr_w_bits_wstrb; // @[BFS.scala 228:12]
  assign io_gather_in_ready = ~vertex_update_buffer_full; // @[BFS.scala 215:54]
  assign io_end = update_engine_io_end; // @[BFS.scala 230:10]
  assign vertex_update_buffer_din = {io_gather_in_bits_tdata,io_level}; // @[Cat.scala 30:58]
  assign vertex_update_buffer_wr_en = io_gather_in_valid & ~FIN; // @[BFS.scala 212:55]
  assign vertex_update_buffer_rd_en = update_engine_io_xbar_in_ready; // @[BFS.scala 225:33]
  assign vertex_update_buffer_clk = clock; // @[BFS.scala 210:46]
  assign vertex_update_buffer_srst = reset; // @[BFS.scala 211:47]
  assign update_engine_clock = clock;
  assign update_engine_reset = reset;
  assign update_engine_io_ddr_aw_ready = io_ddr_aw_ready; // @[BFS.scala 227:13]
  assign update_engine_io_ddr_w_ready = io_ddr_w_ready; // @[BFS.scala 228:12]
  assign update_engine_io_xbar_in_valid = vertex_update_buffer_valid; // @[BFS.scala 219:34]
  assign update_engine_io_xbar_in_bits_tdata = vertex_update_buffer_dout[63:32]; // @[BFS.scala 218:70]
  assign update_engine_io_level_base_addr = io_level_base_addr; // @[BFS.scala 220:36]
  assign update_engine_io_level = vertex_update_buffer_dout[31:0]; // @[BFS.scala 224:57]
  assign update_engine_io_flush = io_flush & _update_engine_io_flush_T; // @[BFS.scala 231:38]
endmodule
module readEdge_engine(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_rdata,
  input  [5:0]   io_in_bits_rid,
  input          io_in_bits_rlast,
  input          io_out_ready,
  output         io_out_valid,
  output [63:0]  io_out_bits_araddr,
  output [5:0]   io_out_bits_arid,
  output [7:0]   io_out_bits_arlen,
  output [2:0]   io_out_bits_arsize,
  input  [63:0]  io_edge_base_addr,
  input  [4:0]   io_free_ptr,
  output [31:0]  io_read_edge_num,
  output         io_read_edge_fifo_empty,
  input  [63:0]  io_inflight_vtxs
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  edge_read_buffer_full; // @[BFS.scala 373:32]
  wire [63:0] edge_read_buffer_din; // @[BFS.scala 373:32]
  wire  edge_read_buffer_wr_en; // @[BFS.scala 373:32]
  wire  edge_read_buffer_empty; // @[BFS.scala 373:32]
  wire [63:0] edge_read_buffer_dout; // @[BFS.scala 373:32]
  wire  edge_read_buffer_rd_en; // @[BFS.scala 373:32]
  wire [5:0] edge_read_buffer_data_count; // @[BFS.scala 373:32]
  wire  edge_read_buffer_clk; // @[BFS.scala 373:32]
  wire  edge_read_buffer_srst; // @[BFS.scala 373:32]
  wire  edge_read_buffer_valid; // @[BFS.scala 373:32]
  reg  transaction_start; // @[BFS.scala 374:34]
  wire  _T = io_in_valid & io_in_ready; // @[BFS.scala 375:20]
  wire  _GEN_0 = _T & io_in_bits_rlast ? 1'h0 : transaction_start; // @[BFS.scala 377:70 BFS.scala 378:23 BFS.scala 374:34]
  wire  _GEN_1 = io_in_valid & io_in_ready & ~io_in_bits_rlast | _GEN_0; // @[BFS.scala 375:66 BFS.scala 376:23]
  wire  _edge_read_buffer_io_wr_en_T_5 = io_in_bits_rdata[63:32] > 32'he; // @[BFS.scala 384:39]
  wire  _edge_read_buffer_io_wr_en_T_6 = ~io_in_bits_rid[5] & io_in_valid & _edge_read_buffer_io_wr_en_T_5; // @[BFS.scala 383:72]
  wire [31:0] remainning_edges = edge_read_buffer_dout[63:32] - 32'he; // @[BFS.scala 388:68]
  reg  cache_status; // @[BFS.scala 393:29]
  reg [31:0] counter; // @[BFS.scala 394:24]
  reg [63:0] araddr; // @[BFS.scala 396:23]
  wire [31:0] next_counter = counter - 32'h40; // @[BFS.scala 398:27]
  wire  _T_10 = ~cache_status; // @[BFS.scala 399:116]
  wire [31:0] _counter_T_1 = remainning_edges - 32'h40; // @[BFS.scala 401:33]
  wire [33:0] _araddr_T_1 = {edge_read_buffer_dout[31:0], 2'h0}; // @[BFS.scala 402:83]
  wire [63:0] _GEN_11 = {{30'd0}, _araddr_T_1}; // @[BFS.scala 402:33]
  wire [63:0] _araddr_T_3 = io_edge_base_addr + _GEN_11; // @[BFS.scala 402:33]
  wire [63:0] _araddr_T_6 = _araddr_T_3 + 64'h100; // @[BFS.scala 402:98]
  wire  _T_15 = counter <= 32'h40; // @[BFS.scala 404:18]
  wire [63:0] _araddr_T_9 = araddr + 64'h100; // @[BFS.scala 410:24]
  wire  _GEN_2 = counter <= 32'h40 ? 1'h0 : cache_status; // @[BFS.scala 404:53 BFS.scala 405:20 BFS.scala 393:29]
  wire  _GEN_5 = io_out_ready & io_out_valid & cache_status ? _GEN_2 : cache_status; // @[BFS.scala 403:82 BFS.scala 393:29]
  wire  _GEN_8 = remainning_edges > 32'h40 & io_out_ready & io_out_valid & ~cache_status | _GEN_5; // @[BFS.scala 399:135 BFS.scala 400:18]
  wire  _num_vertex_T_2 = _T_10 & remainning_edges <= 32'h40; // @[BFS.scala 415:38]
  wire  _num_vertex_T_5 = cache_status & _T_15; // @[BFS.scala 416:42]
  wire [31:0] _num_vertex_T_6 = _num_vertex_T_5 ? counter : 32'h40; // @[Mux.scala 98:16]
  wire [31:0] num_vertex = _num_vertex_T_2 ? remainning_edges : _num_vertex_T_6; // @[Mux.scala 98:16]
  wire [31:0] _arlen_T_1 = {num_vertex[31:2], 2'h0}; // @[BFS.scala 418:63]
  wire [29:0] _arlen_T_6 = num_vertex[31:2] - 30'h1; // @[BFS.scala 420:57]
  wire [29:0] arlen = _arlen_T_1 < num_vertex ? num_vertex[31:2] : _arlen_T_6; // @[BFS.scala 418:18]
  wire  _io_out_valid_T_1 = _T_10 ? edge_read_buffer_valid : 1'h1; // @[BFS.scala 424:22]
  wire  _io_out_valid_T_2 = io_inflight_vtxs < 64'h20; // @[BFS.scala 424:113]
  wire  _io_out_bits_arsize_T = num_vertex <= 32'h1; // @[BFS.scala 429:23]
  wire  _io_out_bits_arsize_T_1 = num_vertex <= 32'h2; // @[BFS.scala 429:23]
  wire [2:0] _io_out_bits_arsize_T_2 = _io_out_bits_arsize_T_1 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  meta_fifo edge_read_buffer ( // @[BFS.scala 373:32]
    .full(edge_read_buffer_full),
    .din(edge_read_buffer_din),
    .wr_en(edge_read_buffer_wr_en),
    .empty(edge_read_buffer_empty),
    .dout(edge_read_buffer_dout),
    .rd_en(edge_read_buffer_rd_en),
    .data_count(edge_read_buffer_data_count),
    .clk(edge_read_buffer_clk),
    .srst(edge_read_buffer_srst),
    .valid(edge_read_buffer_valid)
  );
  assign io_in_ready = ~edge_read_buffer_full; // @[BFS.scala 385:43]
  assign io_out_valid = _io_out_valid_T_1 & io_inflight_vtxs < 64'h20; // @[BFS.scala 424:93]
  assign io_out_bits_araddr = _T_10 ? _araddr_T_3 : araddr; // @[BFS.scala 421:28]
  assign io_out_bits_arid = {1'h1,io_free_ptr}; // @[Cat.scala 30:58]
  assign io_out_bits_arlen = arlen[7:0]; // @[BFS.scala 425:21]
  assign io_out_bits_arsize = _io_out_bits_arsize_T ? 3'h2 : _io_out_bits_arsize_T_2; // @[Mux.scala 98:16]
  assign io_read_edge_num = _num_vertex_T_2 ? remainning_edges : _num_vertex_T_6; // @[Mux.scala 98:16]
  assign io_read_edge_fifo_empty = edge_read_buffer_data_count == 6'h0; // @[util.scala 211:19]
  assign edge_read_buffer_din = io_in_bits_rdata[63:0]; // @[BFS.scala 382:46]
  assign edge_read_buffer_wr_en = _edge_read_buffer_io_wr_en_T_6 & ~transaction_start; // @[BFS.scala 384:61]
  assign edge_read_buffer_rd_en = io_out_ready & _T_10 & _io_out_valid_T_2; // @[BFS.scala 433:79]
  assign edge_read_buffer_clk = clock; // @[BFS.scala 380:42]
  assign edge_read_buffer_srst = reset; // @[BFS.scala 381:43]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 374:34]
      transaction_start <= 1'h0; // @[BFS.scala 374:34]
    end else begin
      transaction_start <= _GEN_1;
    end
    if (reset) begin // @[BFS.scala 393:29]
      cache_status <= 1'h0; // @[BFS.scala 393:29]
    end else begin
      cache_status <= _GEN_8;
    end
    if (reset) begin // @[BFS.scala 394:24]
      counter <= 32'h0; // @[BFS.scala 394:24]
    end else if (remainning_edges > 32'h40 & io_out_ready & io_out_valid & ~cache_status) begin // @[BFS.scala 399:135]
      counter <= _counter_T_1; // @[BFS.scala 401:13]
    end else if (io_out_ready & io_out_valid & cache_status) begin // @[BFS.scala 403:82]
      if (counter <= 32'h40) begin // @[BFS.scala 404:53]
        counter <= 32'h0; // @[BFS.scala 406:15]
      end else begin
        counter <= next_counter; // @[BFS.scala 409:15]
      end
    end
    if (reset) begin // @[BFS.scala 396:23]
      araddr <= 64'h0; // @[BFS.scala 396:23]
    end else if (remainning_edges > 32'h40 & io_out_ready & io_out_valid & ~cache_status) begin // @[BFS.scala 399:135]
      araddr <= _araddr_T_6; // @[BFS.scala 402:12]
    end else if (io_out_ready & io_out_valid & cache_status) begin // @[BFS.scala 403:82]
      if (counter <= 32'h40) begin // @[BFS.scala 404:53]
        araddr <= 64'h0; // @[BFS.scala 407:14]
      end else begin
        araddr <= _araddr_T_9; // @[BFS.scala 410:14]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  transaction_start = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cache_status = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  araddr = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AMBA_Arbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_araddr,
  input  [5:0]  io_in_0_bits_arid,
  input  [7:0]  io_in_0_bits_arlen,
  input  [2:0]  io_in_0_bits_arsize,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_araddr,
  input  [5:0]  io_in_1_bits_arid,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_araddr,
  output [5:0]  io_out_bits_arid,
  output [7:0]  io_out_bits_arlen,
  output [2:0]  io_out_bits_arsize
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  status; // @[util.scala 323:23]
  wire  grant_1 = ~io_in_0_valid; // @[util.scala 312:78]
  reg  grant_reg_0; // @[util.scala 325:26]
  reg  grant_reg_1; // @[util.scala 325:26]
  wire  _T = ~status; // @[util.scala 330:17]
  wire [2:0] _GEN_3 = io_in_0_valid ? io_in_0_bits_arsize : 3'h4; // @[util.scala 331:28 util.scala 333:21 util.scala 328:15]
  wire [7:0] _GEN_4 = io_in_0_valid ? io_in_0_bits_arlen : 8'h3; // @[util.scala 331:28 util.scala 333:21 util.scala 328:15]
  wire [5:0] _GEN_5 = io_in_0_valid ? io_in_0_bits_arid : io_in_1_bits_arid; // @[util.scala 331:28 util.scala 333:21 util.scala 328:15]
  wire [63:0] _GEN_6 = io_in_0_valid ? io_in_0_bits_araddr : io_in_1_bits_araddr; // @[util.scala 331:28 util.scala 333:21 util.scala 328:15]
  wire [2:0] _GEN_10 = grant_reg_0 ? io_in_0_bits_arsize : 3'h4; // @[util.scala 336:26 util.scala 338:21 util.scala 328:15]
  wire [7:0] _GEN_11 = grant_reg_0 ? io_in_0_bits_arlen : 8'h3; // @[util.scala 336:26 util.scala 338:21 util.scala 328:15]
  wire [5:0] _GEN_12 = grant_reg_0 ? io_in_0_bits_arid : io_in_1_bits_arid; // @[util.scala 336:26 util.scala 338:21 util.scala 328:15]
  wire [63:0] _GEN_13 = grant_reg_0 ? io_in_0_bits_araddr : io_in_1_bits_araddr; // @[util.scala 336:26 util.scala 338:21 util.scala 328:15]
  wire [2:0] _GEN_17 = status ? _GEN_10 : 3'h4; // @[util.scala 335:35 util.scala 328:15]
  wire [7:0] _GEN_18 = status ? _GEN_11 : 8'h3; // @[util.scala 335:35 util.scala 328:15]
  wire [5:0] _GEN_19 = status ? _GEN_12 : io_in_1_bits_arid; // @[util.scala 335:35 util.scala 328:15]
  wire [63:0] _GEN_20 = status ? _GEN_13 : io_in_1_bits_araddr; // @[util.scala 335:35 util.scala 328:15]
  wire  _T_8 = grant_1 & io_in_1_valid; // @[util.scala 345:24]
  wire  _GEN_28 = io_out_valid & io_out_ready & status ? 1'h0 : status; // @[util.scala 348:66 util.scala 349:12 util.scala 323:23]
  wire  _GEN_31 = (io_in_0_valid | io_in_1_valid) & _T & ~io_out_ready | _GEN_28; // @[util.scala 343:90 util.scala 347:12]
  assign io_in_0_ready = _T ? io_out_ready : grant_reg_0 & io_out_ready; // @[util.scala 352:20]
  assign io_in_1_ready = _T ? grant_1 & io_out_ready : grant_reg_1 & io_out_ready; // @[util.scala 352:20]
  assign io_out_valid = _T ? ~grant_1 | io_in_1_valid : ~grant_reg_1 | io_in_1_valid; // @[util.scala 354:22]
  assign io_out_bits_araddr = ~status ? _GEN_6 : _GEN_20; // @[util.scala 330:30]
  assign io_out_bits_arid = ~status ? _GEN_5 : _GEN_19; // @[util.scala 330:30]
  assign io_out_bits_arlen = ~status ? _GEN_4 : _GEN_18; // @[util.scala 330:30]
  assign io_out_bits_arsize = ~status ? _GEN_3 : _GEN_17; // @[util.scala 330:30]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 323:23]
      status <= 1'h0; // @[util.scala 323:23]
    end else begin
      status <= _GEN_31;
    end
    if (reset) begin // @[util.scala 325:26]
      grant_reg_0 <= 1'h0; // @[util.scala 325:26]
    end else if ((io_in_0_valid | io_in_1_valid) & _T & ~io_out_ready) begin // @[util.scala 343:90]
      grant_reg_0 <= io_in_0_valid; // @[util.scala 344:15]
    end
    if (reset) begin // @[util.scala 325:26]
      grant_reg_1 <= 1'h0; // @[util.scala 325:26]
    end else if ((io_in_0_valid | io_in_1_valid) & _T & ~io_out_ready) begin // @[util.scala 343:90]
      grant_reg_1 <= _T_8; // @[util.scala 344:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  status = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  grant_reg_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  grant_reg_1 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module regFile(
  input         clock,
  input         reset,
  input  [31:0] io_dataIn,
  output [31:0] io_dataOut,
  input         io_writeFlag,
  input  [4:0]  io_rptr,
  input  [4:0]  io_wptr,
  output [4:0]  io_wcount
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[util.scala 178:21]
  reg [31:0] regs_1; // @[util.scala 178:21]
  reg [31:0] regs_2; // @[util.scala 178:21]
  reg [31:0] regs_3; // @[util.scala 178:21]
  reg [31:0] regs_4; // @[util.scala 178:21]
  reg [31:0] regs_5; // @[util.scala 178:21]
  reg [31:0] regs_6; // @[util.scala 178:21]
  reg [31:0] regs_7; // @[util.scala 178:21]
  reg [31:0] regs_8; // @[util.scala 178:21]
  reg [31:0] regs_9; // @[util.scala 178:21]
  reg [31:0] regs_10; // @[util.scala 178:21]
  reg [31:0] regs_11; // @[util.scala 178:21]
  reg [31:0] regs_12; // @[util.scala 178:21]
  reg [31:0] regs_13; // @[util.scala 178:21]
  reg [31:0] regs_14; // @[util.scala 178:21]
  reg [31:0] regs_15; // @[util.scala 178:21]
  reg [31:0] regs_16; // @[util.scala 178:21]
  reg [31:0] regs_17; // @[util.scala 178:21]
  reg [31:0] regs_18; // @[util.scala 178:21]
  reg [31:0] regs_19; // @[util.scala 178:21]
  reg [31:0] regs_20; // @[util.scala 178:21]
  reg [31:0] regs_21; // @[util.scala 178:21]
  reg [31:0] regs_22; // @[util.scala 178:21]
  reg [31:0] regs_23; // @[util.scala 178:21]
  reg [31:0] regs_24; // @[util.scala 178:21]
  reg [31:0] regs_25; // @[util.scala 178:21]
  reg [31:0] regs_26; // @[util.scala 178:21]
  reg [31:0] regs_27; // @[util.scala 178:21]
  reg [31:0] regs_28; // @[util.scala 178:21]
  reg [31:0] regs_29; // @[util.scala 178:21]
  reg [31:0] regs_30; // @[util.scala 178:21]
  reg [31:0] regs_31; // @[util.scala 178:21]
  wire [31:0] _GEN_1 = 5'h1 == io_rptr ? regs_1 : regs_0; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_2 = 5'h2 == io_rptr ? regs_2 : _GEN_1; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_3 = 5'h3 == io_rptr ? regs_3 : _GEN_2; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_4 = 5'h4 == io_rptr ? regs_4 : _GEN_3; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_5 = 5'h5 == io_rptr ? regs_5 : _GEN_4; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_6 = 5'h6 == io_rptr ? regs_6 : _GEN_5; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_7 = 5'h7 == io_rptr ? regs_7 : _GEN_6; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_8 = 5'h8 == io_rptr ? regs_8 : _GEN_7; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_9 = 5'h9 == io_rptr ? regs_9 : _GEN_8; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_10 = 5'ha == io_rptr ? regs_10 : _GEN_9; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_11 = 5'hb == io_rptr ? regs_11 : _GEN_10; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_12 = 5'hc == io_rptr ? regs_12 : _GEN_11; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_13 = 5'hd == io_rptr ? regs_13 : _GEN_12; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_14 = 5'he == io_rptr ? regs_14 : _GEN_13; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_15 = 5'hf == io_rptr ? regs_15 : _GEN_14; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_16 = 5'h10 == io_rptr ? regs_16 : _GEN_15; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_17 = 5'h11 == io_rptr ? regs_17 : _GEN_16; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_18 = 5'h12 == io_rptr ? regs_18 : _GEN_17; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_19 = 5'h13 == io_rptr ? regs_19 : _GEN_18; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_20 = 5'h14 == io_rptr ? regs_20 : _GEN_19; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_21 = 5'h15 == io_rptr ? regs_21 : _GEN_20; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_22 = 5'h16 == io_rptr ? regs_22 : _GEN_21; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_23 = 5'h17 == io_rptr ? regs_23 : _GEN_22; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_24 = 5'h18 == io_rptr ? regs_24 : _GEN_23; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_25 = 5'h19 == io_rptr ? regs_25 : _GEN_24; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_26 = 5'h1a == io_rptr ? regs_26 : _GEN_25; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_27 = 5'h1b == io_rptr ? regs_27 : _GEN_26; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_28 = 5'h1c == io_rptr ? regs_28 : _GEN_27; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_29 = 5'h1d == io_rptr ? regs_29 : _GEN_28; // @[util.scala 180:14 util.scala 180:14]
  wire [31:0] _GEN_30 = 5'h1e == io_rptr ? regs_30 : _GEN_29; // @[util.scala 180:14 util.scala 180:14]
  reg [4:0] counterValue; // @[Counter.scala 60:40]
  wire [4:0] _wrap_value_T_1 = counterValue + 5'h1; // @[Counter.scala 76:24]
  assign io_dataOut = 5'h1f == io_rptr ? regs_31 : _GEN_30; // @[util.scala 180:14 util.scala 180:14]
  assign io_wcount = counterValue; // @[util.scala 187:13]
  always @(posedge clock) begin
    if (reset) begin // @[util.scala 178:21]
      regs_0 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h0 == io_wptr) begin // @[util.scala 183:19]
        regs_0 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_1 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1 == io_wptr) begin // @[util.scala 183:19]
        regs_1 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_2 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h2 == io_wptr) begin // @[util.scala 183:19]
        regs_2 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_3 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h3 == io_wptr) begin // @[util.scala 183:19]
        regs_3 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_4 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h4 == io_wptr) begin // @[util.scala 183:19]
        regs_4 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_5 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h5 == io_wptr) begin // @[util.scala 183:19]
        regs_5 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_6 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h6 == io_wptr) begin // @[util.scala 183:19]
        regs_6 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_7 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h7 == io_wptr) begin // @[util.scala 183:19]
        regs_7 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_8 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h8 == io_wptr) begin // @[util.scala 183:19]
        regs_8 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_9 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h9 == io_wptr) begin // @[util.scala 183:19]
        regs_9 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_10 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'ha == io_wptr) begin // @[util.scala 183:19]
        regs_10 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_11 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hb == io_wptr) begin // @[util.scala 183:19]
        regs_11 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_12 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hc == io_wptr) begin // @[util.scala 183:19]
        regs_12 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_13 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hd == io_wptr) begin // @[util.scala 183:19]
        regs_13 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_14 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'he == io_wptr) begin // @[util.scala 183:19]
        regs_14 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_15 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'hf == io_wptr) begin // @[util.scala 183:19]
        regs_15 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_16 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h10 == io_wptr) begin // @[util.scala 183:19]
        regs_16 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_17 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h11 == io_wptr) begin // @[util.scala 183:19]
        regs_17 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_18 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h12 == io_wptr) begin // @[util.scala 183:19]
        regs_18 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_19 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h13 == io_wptr) begin // @[util.scala 183:19]
        regs_19 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_20 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h14 == io_wptr) begin // @[util.scala 183:19]
        regs_20 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_21 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h15 == io_wptr) begin // @[util.scala 183:19]
        regs_21 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_22 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h16 == io_wptr) begin // @[util.scala 183:19]
        regs_22 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_23 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h17 == io_wptr) begin // @[util.scala 183:19]
        regs_23 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_24 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h18 == io_wptr) begin // @[util.scala 183:19]
        regs_24 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_25 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h19 == io_wptr) begin // @[util.scala 183:19]
        regs_25 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_26 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1a == io_wptr) begin // @[util.scala 183:19]
        regs_26 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_27 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1b == io_wptr) begin // @[util.scala 183:19]
        regs_27 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_28 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1c == io_wptr) begin // @[util.scala 183:19]
        regs_28 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_29 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1d == io_wptr) begin // @[util.scala 183:19]
        regs_29 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_30 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1e == io_wptr) begin // @[util.scala 183:19]
        regs_30 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[util.scala 178:21]
      regs_31 <= 32'h0; // @[util.scala 178:21]
    end else if (io_writeFlag) begin // @[util.scala 182:21]
      if (5'h1f == io_wptr) begin // @[util.scala 183:19]
        regs_31 <= io_dataIn; // @[util.scala 183:19]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      counterValue <= 5'h0; // @[Counter.scala 60:40]
    end else if (io_writeFlag) begin // @[Counter.scala 118:17]
      counterValue <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  counterValue = _RAND_32[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  input          io_start,
  input  [31:0]  io_root,
  output         io_issue_sync,
  input  [4:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 472:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 472:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 472:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 472:34]
  wire  edge_cache_clock; // @[BFS.scala 481:26]
  wire  edge_cache_reset; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 481:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 481:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 481:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 481:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 481:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 481:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 481:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 481:26]
  wire [4:0] edge_cache_io_free_ptr; // @[BFS.scala 481:26]
  wire [31:0] edge_cache_io_read_edge_num; // @[BFS.scala 481:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_inflight_vtxs; // @[BFS.scala 481:26]
  wire  r_demux_aclk; // @[BFS.scala 485:23]
  wire  r_demux_aresetn; // @[BFS.scala 485:23]
  wire [127:0] r_demux_s_axis_tdata; // @[BFS.scala 485:23]
  wire [15:0] r_demux_s_axis_tkeep; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tlast; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tvalid; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tready; // @[BFS.scala 485:23]
  wire [5:0] r_demux_s_axis_tid; // @[BFS.scala 485:23]
  wire [255:0] r_demux_m_axis_tdata; // @[BFS.scala 485:23]
  wire [31:0] r_demux_m_axis_tkeep; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tlast; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tvalid; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tready; // @[BFS.scala 485:23]
  wire [11:0] r_demux_m_axis_tid; // @[BFS.scala 485:23]
  wire  arbi_clock; // @[BFS.scala 506:20]
  wire  arbi_reset; // @[BFS.scala 506:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 506:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 506:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 506:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 506:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 506:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 506:20]
  wire  arbi_io_out_ready; // @[BFS.scala 506:20]
  wire  arbi_io_out_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 506:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 506:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 506:20]
  wire  num_regfile_clock; // @[BFS.scala 519:27]
  wire  num_regfile_reset; // @[BFS.scala 519:27]
  wire [31:0] num_regfile_io_dataIn; // @[BFS.scala 519:27]
  wire [31:0] num_regfile_io_dataOut; // @[BFS.scala 519:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_wcount; // @[BFS.scala 519:27]
  wire  vertex_out_fifo_full; // @[BFS.scala 581:31]
  wire [131:0] vertex_out_fifo_din; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 581:31]
  wire [131:0] vertex_out_fifo_dout; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 581:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 581:31]
  (*dont_touch = "true" *)reg [2:0] upward_status; // @[BFS.scala 466:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 467:30]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 468:35]
  wire [4:0] vertex_read_id_lo = vertex_read_buffer_data_count[4:0]; // @[BFS.scala 479:76 BFS.scala 479:76]
  wire  r_demux_out_0_valid = r_demux_m_axis_tvalid[0]; // @[BFS.scala 497:42]
  wire [5:0] r_demux_out_0_bits_rid = r_demux_m_axis_tid[5:0]; // @[BFS.scala 498:42]
  wire  r_demux_out_0_bits_rlast = r_demux_m_axis_tlast[0]; // @[BFS.scala 499:46]
  wire [127:0] r_demux_out_0_bits_rdata = r_demux_m_axis_tdata[127:0]; // @[BFS.scala 500:46]
  wire  r_demux_out_1_ready = edge_cache_io_in_ready; // @[BFS.scala 486:25 BFS.scala 504:20]
  wire  r_demux_out_0_ready = ~vertex_out_fifo_full; // @[BFS.scala 594:51]
  wire [37:0] _arbi_io_in_1_bits_araddr_T = {vertex_read_buffer_dout, 6'h0}; // @[BFS.scala 508:86]
  wire [63:0] _GEN_31 = {{26'd0}, _arbi_io_in_1_bits_araddr_T}; // @[BFS.scala 508:56]
  wire  _arbi_io_in_1_valid_T_3 = inflight_vtxs < 64'h20; // @[BFS.scala 509:116]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 515:96]
  reg [1:0] status; // @[BFS.scala 534:23]
  reg [31:0] num; // @[BFS.scala 535:20]
  wire  _T = status == 2'h0; // @[BFS.scala 536:15]
  wire  _T_4 = status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready; // @[BFS.scala 536:66]
  wire  _T_8 = status == 2'h2; // @[BFS.scala 544:22]
  wire  _T_9 = status == 2'h1; // @[BFS.scala 544:60]
  wire  _T_10 = status == 2'h2 | status == 2'h1; // @[BFS.scala 544:50]
  wire [31:0] _num_T_2 = num - 32'h4; // @[BFS.scala 560:18]
  wire [31:0] _num_T_6 = num > 32'h4 ? _num_T_2 : 32'h0; // @[BFS.scala 566:17]
  wire [31:0] _GEN_6 = r_demux_out_0_bits_rlast ? 32'h0 : _num_T_6; // @[BFS.scala 563:45 BFS.scala 564:11 BFS.scala 566:11]
  wire  _keep_0_T_3 = _T & r_demux_out_0_bits_rid[5]; // @[BFS.scala 573:33]
  wire  _keep_0_T_4 = num_regfile_io_dataOut > 32'h0; // @[BFS.scala 573:109]
  wire  _keep_0_T_6 = num > 32'h0; // @[BFS.scala 574:51]
  wire  _keep_0_T_10 = ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 575:36]
  wire  _keep_0_T_11 = _T & ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 575:33]
  wire [31:0] _keep_0_T_15 = r_demux_out_0_bits_rdata[63:32] + 32'h2; // @[BFS.scala 576:80]
  wire [2:0] _keep_0_T_22 = 3'h4 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_32 = {{29'd0}, _keep_0_T_22}; // @[BFS.scala 577:56]
  wire  _keep_0_T_23 = num > _GEN_32; // @[BFS.scala 577:56]
  wire  _keep_0_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_0_T_23; // @[Mux.scala 98:16]
  wire  _keep_0_T_26 = _T_8 ? _keep_0_T_6 : _keep_0_T_25; // @[Mux.scala 98:16]
  wire  keep_0 = _keep_0_T_3 ? _keep_0_T_4 : _keep_0_T_26; // @[Mux.scala 98:16]
  wire  _keep_1_T_4 = num_regfile_io_dataOut > 32'h1; // @[BFS.scala 573:109]
  wire  _keep_1_T_6 = num > 32'h1; // @[BFS.scala 574:51]
  wire [2:0] _keep_1_T_22 = 3'h5 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_33 = {{29'd0}, _keep_1_T_22}; // @[BFS.scala 577:56]
  wire  _keep_1_T_23 = num > _GEN_33; // @[BFS.scala 577:56]
  wire  _keep_1_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_1_T_23; // @[Mux.scala 98:16]
  wire  _keep_1_T_26 = _T_8 ? _keep_1_T_6 : _keep_1_T_25; // @[Mux.scala 98:16]
  wire  keep_1 = _keep_0_T_3 ? _keep_1_T_4 : _keep_1_T_26; // @[Mux.scala 98:16]
  wire  _keep_2_T_4 = num_regfile_io_dataOut > 32'h2; // @[BFS.scala 573:109]
  wire  _keep_2_T_6 = num > 32'h2; // @[BFS.scala 574:51]
  wire  _keep_2_T_16 = _keep_0_T_15 > 32'h2; // @[BFS.scala 576:87]
  wire [2:0] _keep_2_T_22 = 3'h6 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_34 = {{29'd0}, _keep_2_T_22}; // @[BFS.scala 577:56]
  wire  _keep_2_T_23 = num > _GEN_34; // @[BFS.scala 577:56]
  wire  _keep_2_T_25 = _keep_0_T_11 ? _keep_2_T_16 : _T_9 & _keep_2_T_23; // @[Mux.scala 98:16]
  wire  _keep_2_T_26 = _T_8 ? _keep_2_T_6 : _keep_2_T_25; // @[Mux.scala 98:16]
  wire  keep_2 = _keep_0_T_3 ? _keep_2_T_4 : _keep_2_T_26; // @[Mux.scala 98:16]
  wire  _keep_3_T_4 = num_regfile_io_dataOut > 32'h3; // @[BFS.scala 573:109]
  wire  _keep_3_T_6 = num > 32'h3; // @[BFS.scala 574:51]
  wire  _keep_3_T_16 = _keep_0_T_15 > 32'h3; // @[BFS.scala 576:87]
  wire [2:0] _keep_3_T_22 = 3'h7 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_35 = {{29'd0}, _keep_3_T_22}; // @[BFS.scala 577:56]
  wire  _keep_3_T_23 = num > _GEN_35; // @[BFS.scala 577:56]
  wire  _keep_3_T_25 = _keep_0_T_11 ? _keep_3_T_16 : _T_9 & _keep_3_T_23; // @[Mux.scala 98:16]
  wire  _keep_3_T_26 = _T_8 ? _keep_3_T_6 : _keep_3_T_25; // @[Mux.scala 98:16]
  wire  keep_3 = _keep_0_T_3 ? _keep_3_T_4 : _keep_3_T_26; // @[Mux.scala 98:16]
  wire [131:0] _vertex_out_fifo_io_din_T = {r_demux_out_0_bits_rdata,keep_3,keep_2,keep_1,keep_0}; // @[Cat.scala 30:58]
  wire [35:0] _vertex_out_fifo_io_din_T_1 = {io_root,4'h1}; // @[Cat.scala 30:58]
  wire [131:0] _vertex_out_fifo_io_din_T_4 = _vertex_read_buffer_io_rd_en_T_2 ? 132'h800000001 :
    _vertex_out_fifo_io_din_T; // @[Mux.scala 98:16]
  reg  syncRecv_0; // @[BFS.scala 597:25]
  reg  syncRecv_1; // @[BFS.scala 597:25]
  reg  syncRecv_2; // @[BFS.scala 597:25]
  reg  syncRecv_3; // @[BFS.scala 597:25]
  reg  syncRecv_4; // @[BFS.scala 597:25]
  wire  _GEN_10 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_12 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_14 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_16 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_18 = io_recv_sync[4] | syncRecv_4; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 607:34]
  wire [31:0] _T_47 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_51 = _T_47[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_61 = vertex_out_fifo_data_count == 6'h0; // @[util.scala 211:19]
  wire  _T_62 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_61; // @[BFS.scala 612:71]
  wire [2:0] _GEN_21 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 621:53 BFS.scala 622:19 BFS.scala 466:30]
  wire [2:0] _GEN_22 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3 & syncRecv_4) ? 3'h3 :
    _GEN_21; // @[BFS.scala 615:71]
  wire  _T_79 = r_demux_out_0_valid & r_demux_out_0_ready & _keep_0_T_10; // @[BFS.scala 627:77]
  wire [63:0] _GEN_37 = {{32'd0}, r_demux_out_0_bits_rdata[63:32]}; // @[BFS.scala 629:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_37; // @[BFS.scala 629:46]
  wire  _T_82 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 632:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 636:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 638:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 472:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 481:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_free_ptr(edge_cache_io_free_ptr),
    .io_read_edge_num(edge_cache_io_read_edge_num),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_inflight_vtxs(edge_cache_io_inflight_vtxs)
  );
  r_demux r_demux ( // @[BFS.scala 485:23]
    .aclk(r_demux_aclk),
    .aresetn(r_demux_aresetn),
    .s_axis_tdata(r_demux_s_axis_tdata),
    .s_axis_tkeep(r_demux_s_axis_tkeep),
    .s_axis_tlast(r_demux_s_axis_tlast),
    .s_axis_tvalid(r_demux_s_axis_tvalid),
    .s_axis_tready(r_demux_s_axis_tready),
    .s_axis_tid(r_demux_s_axis_tid),
    .m_axis_tdata(r_demux_m_axis_tdata),
    .m_axis_tkeep(r_demux_m_axis_tkeep),
    .m_axis_tlast(r_demux_m_axis_tlast),
    .m_axis_tvalid(r_demux_m_axis_tvalid),
    .m_axis_tready(r_demux_m_axis_tready),
    .m_axis_tid(r_demux_m_axis_tid)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 506:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  regFile num_regfile ( // @[BFS.scala 519:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr),
    .io_wcount(num_regfile_io_wcount)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 581:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 507:13]
  assign io_ddr_r_ready = r_demux_s_axis_tready; // @[BFS.scala 494:18]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 477:52]
  assign io_xbar_out_valid = vertex_out_fifo_valid; // @[BFS.scala 584:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_dout[131:4]; // @[BFS.scala 586:52]
  assign io_xbar_out_bits_tkeep = vertex_out_fifo_dout[3:0]; // @[BFS.scala 585:52]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 469:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 607:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 476:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 475:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 515:80]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 473:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 474:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = r_demux_m_axis_tvalid[1]; // @[BFS.scala 497:42]
  assign edge_cache_io_in_bits_rdata = r_demux_m_axis_tdata[255:128]; // @[BFS.scala 500:46]
  assign edge_cache_io_in_bits_rid = r_demux_m_axis_tid[11:6]; // @[BFS.scala 498:42]
  assign edge_cache_io_in_bits_rlast = r_demux_m_axis_tlast[1]; // @[BFS.scala 499:46]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 516:17]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 483:32]
  assign edge_cache_io_free_ptr = num_regfile_io_wcount; // @[BFS.scala 524:26]
  assign edge_cache_io_inflight_vtxs = inflight_vtxs; // @[BFS.scala 484:31]
  assign r_demux_aclk = clock; // @[BFS.scala 492:34]
  assign r_demux_aresetn = ~reset; // @[BFS.scala 493:25]
  assign r_demux_s_axis_tdata = io_ddr_r_bits_rdata; // @[BFS.scala 488:27]
  assign r_demux_s_axis_tkeep = 16'hffff; // @[nf_arm_doce_top.scala 128:85]
  assign r_demux_s_axis_tlast = io_ddr_r_bits_rlast; // @[BFS.scala 489:27]
  assign r_demux_s_axis_tvalid = io_ddr_r_valid; // @[BFS.scala 487:28]
  assign r_demux_s_axis_tid = io_ddr_r_bits_rid; // @[BFS.scala 491:25]
  assign r_demux_m_axis_tready = {r_demux_out_1_ready,r_demux_out_0_ready}; // @[BFS.scala 503:84]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 516:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & inflight_vtxs < 64'h20; // @[BFS.scala 509:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_31; // @[BFS.scala 508:56]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id_lo}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 507:13]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = edge_cache_io_read_edge_num; // @[BFS.scala 522:25]
  assign num_regfile_io_writeFlag = arbi_io_in_0_ready & arbi_io_in_0_valid; // @[BFS.scala 520:51]
  assign num_regfile_io_rptr = r_demux_out_0_bits_rid[4:0]; // @[BFS.scala 369:7]
  assign num_regfile_io_wptr = num_regfile_io_wcount; // @[BFS.scala 521:23]
  assign vertex_out_fifo_din = io_start ? {{96'd0}, _vertex_out_fifo_io_din_T_1} : _vertex_out_fifo_io_din_T_4; // @[Mux.scala 98:16]
  assign vertex_out_fifo_wr_en = r_demux_out_0_valid | _vertex_read_buffer_io_rd_en_T_2 | io_start; // @[BFS.scala 589:93]
  assign vertex_out_fifo_rd_en = io_xbar_out_ready; // @[BFS.scala 588:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 583:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 582:42]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 466:30]
      upward_status <= 3'h0; // @[BFS.scala 466:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 608:57]
      upward_status <= 3'h1; // @[BFS.scala 609:19]
    end else if (upward_status == 3'h1 & (_T_51 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3 | syncRecv_4))
      ) begin // @[BFS.scala 610:105]
      upward_status <= 3'h2; // @[BFS.scala 611:19]
    end else if (_T_62 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 613:62]
      upward_status <= 3'h4; // @[BFS.scala 614:19]
    end else begin
      upward_status <= _GEN_22;
    end
    if (reset) begin // @[BFS.scala 467:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 467:30]
    end else if (!(_T_82 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 633:91]
      if (_T_82) begin // @[BFS.scala 635:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 636:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 637:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 638:19]
      end
    end
    if (reset) begin // @[BFS.scala 468:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 468:35]
    end else if (io_signal) begin // @[BFS.scala 625:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 626:24]
    end else if (_T_79 & _T) begin // @[BFS.scala 628:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 629:24]
    end
    if (reset) begin // @[BFS.scala 534:23]
      status <= 2'h0; // @[BFS.scala 534:23]
    end else if (status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 536:99]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 537:45]
        status <= 2'h0; // @[BFS.scala 538:14]
      end else if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 539:61]
        status <= 2'h2; // @[BFS.scala 540:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 542:14]
      end
    end else if (_T_10 & r_demux_out_0_valid & r_demux_out_0_ready & r_demux_out_0_bits_rlast) begin // @[BFS.scala 545:117]
      status <= 2'h0; // @[BFS.scala 546:14]
    end
    if (reset) begin // @[BFS.scala 535:20]
      num <= 32'h0; // @[BFS.scala 535:20]
    end else if (_T_4 & ~r_demux_out_0_bits_rlast) begin // @[BFS.scala 550:112]
      if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 551:55]
        num <= num_regfile_io_dataOut; // @[BFS.scala 552:11]
      end else begin
        num <= r_demux_out_0_bits_rdata[63:32]; // @[BFS.scala 554:11]
      end
    end else if (_T_8 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 556:114]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 557:45]
        num <= 32'h0; // @[BFS.scala 558:11]
      end else begin
        num <= _num_T_2; // @[BFS.scala 560:11]
      end
    end else if (_T_9 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 562:119]
      num <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_0 <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_1 <= _GEN_12;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_2 <= _GEN_14;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_3 <= _GEN_16;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_4 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_4 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_4 <= _GEN_18;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  status = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  num = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  syncRecv_4 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_1(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [4:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 472:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 472:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 472:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 472:34]
  wire  edge_cache_clock; // @[BFS.scala 481:26]
  wire  edge_cache_reset; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 481:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 481:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 481:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 481:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 481:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 481:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 481:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 481:26]
  wire [4:0] edge_cache_io_free_ptr; // @[BFS.scala 481:26]
  wire [31:0] edge_cache_io_read_edge_num; // @[BFS.scala 481:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_inflight_vtxs; // @[BFS.scala 481:26]
  wire  r_demux_aclk; // @[BFS.scala 485:23]
  wire  r_demux_aresetn; // @[BFS.scala 485:23]
  wire [127:0] r_demux_s_axis_tdata; // @[BFS.scala 485:23]
  wire [15:0] r_demux_s_axis_tkeep; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tlast; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tvalid; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tready; // @[BFS.scala 485:23]
  wire [5:0] r_demux_s_axis_tid; // @[BFS.scala 485:23]
  wire [255:0] r_demux_m_axis_tdata; // @[BFS.scala 485:23]
  wire [31:0] r_demux_m_axis_tkeep; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tlast; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tvalid; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tready; // @[BFS.scala 485:23]
  wire [11:0] r_demux_m_axis_tid; // @[BFS.scala 485:23]
  wire  arbi_clock; // @[BFS.scala 506:20]
  wire  arbi_reset; // @[BFS.scala 506:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 506:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 506:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 506:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 506:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 506:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 506:20]
  wire  arbi_io_out_ready; // @[BFS.scala 506:20]
  wire  arbi_io_out_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 506:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 506:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 506:20]
  wire  num_regfile_clock; // @[BFS.scala 519:27]
  wire  num_regfile_reset; // @[BFS.scala 519:27]
  wire [31:0] num_regfile_io_dataIn; // @[BFS.scala 519:27]
  wire [31:0] num_regfile_io_dataOut; // @[BFS.scala 519:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_wcount; // @[BFS.scala 519:27]
  wire  vertex_out_fifo_full; // @[BFS.scala 581:31]
  wire [131:0] vertex_out_fifo_din; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 581:31]
  wire [131:0] vertex_out_fifo_dout; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 581:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 581:31]
  (*dont_touch = "true" *)reg [2:0] upward_status; // @[BFS.scala 466:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 467:30]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 468:35]
  wire [4:0] vertex_read_id_lo = vertex_read_buffer_data_count[4:0]; // @[BFS.scala 479:76 BFS.scala 479:76]
  wire  r_demux_out_0_valid = r_demux_m_axis_tvalid[0]; // @[BFS.scala 497:42]
  wire [5:0] r_demux_out_0_bits_rid = r_demux_m_axis_tid[5:0]; // @[BFS.scala 498:42]
  wire  r_demux_out_0_bits_rlast = r_demux_m_axis_tlast[0]; // @[BFS.scala 499:46]
  wire [127:0] r_demux_out_0_bits_rdata = r_demux_m_axis_tdata[127:0]; // @[BFS.scala 500:46]
  wire  r_demux_out_1_ready = edge_cache_io_in_ready; // @[BFS.scala 486:25 BFS.scala 504:20]
  wire  r_demux_out_0_ready = ~vertex_out_fifo_full; // @[BFS.scala 594:51]
  wire [37:0] _arbi_io_in_1_bits_araddr_T = {vertex_read_buffer_dout, 6'h0}; // @[BFS.scala 508:86]
  wire [63:0] _GEN_31 = {{26'd0}, _arbi_io_in_1_bits_araddr_T}; // @[BFS.scala 508:56]
  wire  _arbi_io_in_1_valid_T_3 = inflight_vtxs < 64'h20; // @[BFS.scala 509:116]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 515:96]
  reg [1:0] status; // @[BFS.scala 534:23]
  reg [31:0] num; // @[BFS.scala 535:20]
  wire  _T = status == 2'h0; // @[BFS.scala 536:15]
  wire  _T_4 = status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready; // @[BFS.scala 536:66]
  wire  _T_8 = status == 2'h2; // @[BFS.scala 544:22]
  wire  _T_9 = status == 2'h1; // @[BFS.scala 544:60]
  wire  _T_10 = status == 2'h2 | status == 2'h1; // @[BFS.scala 544:50]
  wire [31:0] _num_T_2 = num - 32'h4; // @[BFS.scala 560:18]
  wire [31:0] _num_T_6 = num > 32'h4 ? _num_T_2 : 32'h0; // @[BFS.scala 566:17]
  wire [31:0] _GEN_6 = r_demux_out_0_bits_rlast ? 32'h0 : _num_T_6; // @[BFS.scala 563:45 BFS.scala 564:11 BFS.scala 566:11]
  wire  _keep_0_T_3 = _T & r_demux_out_0_bits_rid[5]; // @[BFS.scala 573:33]
  wire  _keep_0_T_4 = num_regfile_io_dataOut > 32'h0; // @[BFS.scala 573:109]
  wire  _keep_0_T_6 = num > 32'h0; // @[BFS.scala 574:51]
  wire  _keep_0_T_10 = ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 575:36]
  wire  _keep_0_T_11 = _T & ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 575:33]
  wire [31:0] _keep_0_T_15 = r_demux_out_0_bits_rdata[63:32] + 32'h2; // @[BFS.scala 576:80]
  wire [2:0] _keep_0_T_22 = 3'h4 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_32 = {{29'd0}, _keep_0_T_22}; // @[BFS.scala 577:56]
  wire  _keep_0_T_23 = num > _GEN_32; // @[BFS.scala 577:56]
  wire  _keep_0_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_0_T_23; // @[Mux.scala 98:16]
  wire  _keep_0_T_26 = _T_8 ? _keep_0_T_6 : _keep_0_T_25; // @[Mux.scala 98:16]
  wire  keep_0 = _keep_0_T_3 ? _keep_0_T_4 : _keep_0_T_26; // @[Mux.scala 98:16]
  wire  _keep_1_T_4 = num_regfile_io_dataOut > 32'h1; // @[BFS.scala 573:109]
  wire  _keep_1_T_6 = num > 32'h1; // @[BFS.scala 574:51]
  wire [2:0] _keep_1_T_22 = 3'h5 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_33 = {{29'd0}, _keep_1_T_22}; // @[BFS.scala 577:56]
  wire  _keep_1_T_23 = num > _GEN_33; // @[BFS.scala 577:56]
  wire  _keep_1_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_1_T_23; // @[Mux.scala 98:16]
  wire  _keep_1_T_26 = _T_8 ? _keep_1_T_6 : _keep_1_T_25; // @[Mux.scala 98:16]
  wire  keep_1 = _keep_0_T_3 ? _keep_1_T_4 : _keep_1_T_26; // @[Mux.scala 98:16]
  wire  _keep_2_T_4 = num_regfile_io_dataOut > 32'h2; // @[BFS.scala 573:109]
  wire  _keep_2_T_6 = num > 32'h2; // @[BFS.scala 574:51]
  wire  _keep_2_T_16 = _keep_0_T_15 > 32'h2; // @[BFS.scala 576:87]
  wire [2:0] _keep_2_T_22 = 3'h6 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_34 = {{29'd0}, _keep_2_T_22}; // @[BFS.scala 577:56]
  wire  _keep_2_T_23 = num > _GEN_34; // @[BFS.scala 577:56]
  wire  _keep_2_T_25 = _keep_0_T_11 ? _keep_2_T_16 : _T_9 & _keep_2_T_23; // @[Mux.scala 98:16]
  wire  _keep_2_T_26 = _T_8 ? _keep_2_T_6 : _keep_2_T_25; // @[Mux.scala 98:16]
  wire  keep_2 = _keep_0_T_3 ? _keep_2_T_4 : _keep_2_T_26; // @[Mux.scala 98:16]
  wire  _keep_3_T_4 = num_regfile_io_dataOut > 32'h3; // @[BFS.scala 573:109]
  wire  _keep_3_T_6 = num > 32'h3; // @[BFS.scala 574:51]
  wire  _keep_3_T_16 = _keep_0_T_15 > 32'h3; // @[BFS.scala 576:87]
  wire [2:0] _keep_3_T_22 = 3'h7 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_35 = {{29'd0}, _keep_3_T_22}; // @[BFS.scala 577:56]
  wire  _keep_3_T_23 = num > _GEN_35; // @[BFS.scala 577:56]
  wire  _keep_3_T_25 = _keep_0_T_11 ? _keep_3_T_16 : _T_9 & _keep_3_T_23; // @[Mux.scala 98:16]
  wire  _keep_3_T_26 = _T_8 ? _keep_3_T_6 : _keep_3_T_25; // @[Mux.scala 98:16]
  wire  keep_3 = _keep_0_T_3 ? _keep_3_T_4 : _keep_3_T_26; // @[Mux.scala 98:16]
  wire [131:0] _vertex_out_fifo_io_din_T = {r_demux_out_0_bits_rdata,keep_3,keep_2,keep_1,keep_0}; // @[Cat.scala 30:58]
  reg  syncRecv_0; // @[BFS.scala 597:25]
  reg  syncRecv_1; // @[BFS.scala 597:25]
  reg  syncRecv_2; // @[BFS.scala 597:25]
  reg  syncRecv_3; // @[BFS.scala 597:25]
  reg  syncRecv_4; // @[BFS.scala 597:25]
  wire  _GEN_10 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_12 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_14 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_16 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_18 = io_recv_sync[4] | syncRecv_4; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 607:34]
  wire [31:0] _T_47 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_51 = _T_47[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_61 = vertex_out_fifo_data_count == 6'h0; // @[util.scala 211:19]
  wire  _T_62 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_61; // @[BFS.scala 612:71]
  wire [2:0] _GEN_21 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 621:53 BFS.scala 622:19 BFS.scala 466:30]
  wire [2:0] _GEN_22 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3 & syncRecv_4) ? 3'h0 :
    _GEN_21; // @[BFS.scala 615:71]
  wire  _T_79 = r_demux_out_0_valid & r_demux_out_0_ready & _keep_0_T_10; // @[BFS.scala 627:77]
  wire [63:0] _GEN_37 = {{32'd0}, r_demux_out_0_bits_rdata[63:32]}; // @[BFS.scala 629:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_37; // @[BFS.scala 629:46]
  wire  _T_82 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 632:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 636:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 638:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 472:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 481:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_free_ptr(edge_cache_io_free_ptr),
    .io_read_edge_num(edge_cache_io_read_edge_num),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_inflight_vtxs(edge_cache_io_inflight_vtxs)
  );
  r_demux r_demux ( // @[BFS.scala 485:23]
    .aclk(r_demux_aclk),
    .aresetn(r_demux_aresetn),
    .s_axis_tdata(r_demux_s_axis_tdata),
    .s_axis_tkeep(r_demux_s_axis_tkeep),
    .s_axis_tlast(r_demux_s_axis_tlast),
    .s_axis_tvalid(r_demux_s_axis_tvalid),
    .s_axis_tready(r_demux_s_axis_tready),
    .s_axis_tid(r_demux_s_axis_tid),
    .m_axis_tdata(r_demux_m_axis_tdata),
    .m_axis_tkeep(r_demux_m_axis_tkeep),
    .m_axis_tlast(r_demux_m_axis_tlast),
    .m_axis_tvalid(r_demux_m_axis_tvalid),
    .m_axis_tready(r_demux_m_axis_tready),
    .m_axis_tid(r_demux_m_axis_tid)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 506:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  regFile num_regfile ( // @[BFS.scala 519:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr),
    .io_wcount(num_regfile_io_wcount)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 581:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 507:13]
  assign io_ddr_r_ready = r_demux_s_axis_tready; // @[BFS.scala 494:18]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 477:52]
  assign io_xbar_out_valid = vertex_out_fifo_valid; // @[BFS.scala 584:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_dout[131:4]; // @[BFS.scala 586:52]
  assign io_xbar_out_bits_tkeep = vertex_out_fifo_dout[3:0]; // @[BFS.scala 585:52]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 469:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 607:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 476:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 475:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 515:80]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 473:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 474:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = r_demux_m_axis_tvalid[1]; // @[BFS.scala 497:42]
  assign edge_cache_io_in_bits_rdata = r_demux_m_axis_tdata[255:128]; // @[BFS.scala 500:46]
  assign edge_cache_io_in_bits_rid = r_demux_m_axis_tid[11:6]; // @[BFS.scala 498:42]
  assign edge_cache_io_in_bits_rlast = r_demux_m_axis_tlast[1]; // @[BFS.scala 499:46]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 516:17]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 483:32]
  assign edge_cache_io_free_ptr = num_regfile_io_wcount; // @[BFS.scala 524:26]
  assign edge_cache_io_inflight_vtxs = inflight_vtxs; // @[BFS.scala 484:31]
  assign r_demux_aclk = clock; // @[BFS.scala 492:34]
  assign r_demux_aresetn = ~reset; // @[BFS.scala 493:25]
  assign r_demux_s_axis_tdata = io_ddr_r_bits_rdata; // @[BFS.scala 488:27]
  assign r_demux_s_axis_tkeep = 16'hffff; // @[nf_arm_doce_top.scala 128:85]
  assign r_demux_s_axis_tlast = io_ddr_r_bits_rlast; // @[BFS.scala 489:27]
  assign r_demux_s_axis_tvalid = io_ddr_r_valid; // @[BFS.scala 487:28]
  assign r_demux_s_axis_tid = io_ddr_r_bits_rid; // @[BFS.scala 491:25]
  assign r_demux_m_axis_tready = {r_demux_out_1_ready,r_demux_out_0_ready}; // @[BFS.scala 503:84]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 516:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & inflight_vtxs < 64'h20; // @[BFS.scala 509:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_31; // @[BFS.scala 508:56]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id_lo}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 507:13]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = edge_cache_io_read_edge_num; // @[BFS.scala 522:25]
  assign num_regfile_io_writeFlag = arbi_io_in_0_ready & arbi_io_in_0_valid; // @[BFS.scala 520:51]
  assign num_regfile_io_rptr = r_demux_out_0_bits_rid[4:0]; // @[BFS.scala 369:7]
  assign num_regfile_io_wptr = num_regfile_io_wcount; // @[BFS.scala 521:23]
  assign vertex_out_fifo_din = _vertex_read_buffer_io_rd_en_T_2 ? 132'h800000001 : _vertex_out_fifo_io_din_T; // @[Mux.scala 98:16]
  assign vertex_out_fifo_wr_en = r_demux_out_0_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 589:52]
  assign vertex_out_fifo_rd_en = io_xbar_out_ready; // @[BFS.scala 588:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 583:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 582:42]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 466:30]
      upward_status <= 3'h0; // @[BFS.scala 466:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 608:57]
      upward_status <= 3'h1; // @[BFS.scala 609:19]
    end else if (upward_status == 3'h1 & (_T_51 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3 | syncRecv_4))
      ) begin // @[BFS.scala 610:105]
      upward_status <= 3'h2; // @[BFS.scala 611:19]
    end else if (_T_62 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 613:62]
      upward_status <= 3'h4; // @[BFS.scala 614:19]
    end else begin
      upward_status <= _GEN_22;
    end
    if (reset) begin // @[BFS.scala 467:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 467:30]
    end else if (!(_T_82 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 633:91]
      if (_T_82) begin // @[BFS.scala 635:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 636:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 637:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 638:19]
      end
    end
    if (reset) begin // @[BFS.scala 468:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 468:35]
    end else if (io_signal) begin // @[BFS.scala 625:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 626:24]
    end else if (_T_79 & _T) begin // @[BFS.scala 628:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 629:24]
    end
    if (reset) begin // @[BFS.scala 534:23]
      status <= 2'h0; // @[BFS.scala 534:23]
    end else if (status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 536:99]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 537:45]
        status <= 2'h0; // @[BFS.scala 538:14]
      end else if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 539:61]
        status <= 2'h2; // @[BFS.scala 540:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 542:14]
      end
    end else if (_T_10 & r_demux_out_0_valid & r_demux_out_0_ready & r_demux_out_0_bits_rlast) begin // @[BFS.scala 545:117]
      status <= 2'h0; // @[BFS.scala 546:14]
    end
    if (reset) begin // @[BFS.scala 535:20]
      num <= 32'h0; // @[BFS.scala 535:20]
    end else if (_T_4 & ~r_demux_out_0_bits_rlast) begin // @[BFS.scala 550:112]
      if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 551:55]
        num <= num_regfile_io_dataOut; // @[BFS.scala 552:11]
      end else begin
        num <= r_demux_out_0_bits_rdata[63:32]; // @[BFS.scala 554:11]
      end
    end else if (_T_8 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 556:114]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 557:45]
        num <= 32'h0; // @[BFS.scala 558:11]
      end else begin
        num <= _num_T_2; // @[BFS.scala 560:11]
      end
    end else if (_T_9 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 562:119]
      num <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_0 <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_1 <= _GEN_12;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_2 <= _GEN_14;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_3 <= _GEN_16;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_4 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_4 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_4 <= _GEN_18;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  status = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  num = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  syncRecv_4 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_2(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [4:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 472:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 472:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 472:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 472:34]
  wire  edge_cache_clock; // @[BFS.scala 481:26]
  wire  edge_cache_reset; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 481:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 481:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 481:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 481:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 481:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 481:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 481:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 481:26]
  wire [4:0] edge_cache_io_free_ptr; // @[BFS.scala 481:26]
  wire [31:0] edge_cache_io_read_edge_num; // @[BFS.scala 481:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_inflight_vtxs; // @[BFS.scala 481:26]
  wire  r_demux_aclk; // @[BFS.scala 485:23]
  wire  r_demux_aresetn; // @[BFS.scala 485:23]
  wire [127:0] r_demux_s_axis_tdata; // @[BFS.scala 485:23]
  wire [15:0] r_demux_s_axis_tkeep; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tlast; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tvalid; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tready; // @[BFS.scala 485:23]
  wire [5:0] r_demux_s_axis_tid; // @[BFS.scala 485:23]
  wire [255:0] r_demux_m_axis_tdata; // @[BFS.scala 485:23]
  wire [31:0] r_demux_m_axis_tkeep; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tlast; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tvalid; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tready; // @[BFS.scala 485:23]
  wire [11:0] r_demux_m_axis_tid; // @[BFS.scala 485:23]
  wire  arbi_clock; // @[BFS.scala 506:20]
  wire  arbi_reset; // @[BFS.scala 506:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 506:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 506:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 506:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 506:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 506:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 506:20]
  wire  arbi_io_out_ready; // @[BFS.scala 506:20]
  wire  arbi_io_out_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 506:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 506:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 506:20]
  wire  num_regfile_clock; // @[BFS.scala 519:27]
  wire  num_regfile_reset; // @[BFS.scala 519:27]
  wire [31:0] num_regfile_io_dataIn; // @[BFS.scala 519:27]
  wire [31:0] num_regfile_io_dataOut; // @[BFS.scala 519:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_wcount; // @[BFS.scala 519:27]
  wire  vertex_out_fifo_full; // @[BFS.scala 581:31]
  wire [131:0] vertex_out_fifo_din; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 581:31]
  wire [131:0] vertex_out_fifo_dout; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 581:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 581:31]
  (*dont_touch = "true" *)reg [2:0] upward_status; // @[BFS.scala 466:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 467:30]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 468:35]
  wire [4:0] vertex_read_id_lo = vertex_read_buffer_data_count[4:0]; // @[BFS.scala 479:76 BFS.scala 479:76]
  wire  r_demux_out_0_valid = r_demux_m_axis_tvalid[0]; // @[BFS.scala 497:42]
  wire [5:0] r_demux_out_0_bits_rid = r_demux_m_axis_tid[5:0]; // @[BFS.scala 498:42]
  wire  r_demux_out_0_bits_rlast = r_demux_m_axis_tlast[0]; // @[BFS.scala 499:46]
  wire [127:0] r_demux_out_0_bits_rdata = r_demux_m_axis_tdata[127:0]; // @[BFS.scala 500:46]
  wire  r_demux_out_1_ready = edge_cache_io_in_ready; // @[BFS.scala 486:25 BFS.scala 504:20]
  wire  r_demux_out_0_ready = ~vertex_out_fifo_full; // @[BFS.scala 594:51]
  wire [37:0] _arbi_io_in_1_bits_araddr_T = {vertex_read_buffer_dout, 6'h0}; // @[BFS.scala 508:86]
  wire [63:0] _GEN_31 = {{26'd0}, _arbi_io_in_1_bits_araddr_T}; // @[BFS.scala 508:56]
  wire  _arbi_io_in_1_valid_T_3 = inflight_vtxs < 64'h20; // @[BFS.scala 509:116]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 515:96]
  reg [1:0] status; // @[BFS.scala 534:23]
  reg [31:0] num; // @[BFS.scala 535:20]
  wire  _T = status == 2'h0; // @[BFS.scala 536:15]
  wire  _T_4 = status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready; // @[BFS.scala 536:66]
  wire  _T_8 = status == 2'h2; // @[BFS.scala 544:22]
  wire  _T_9 = status == 2'h1; // @[BFS.scala 544:60]
  wire  _T_10 = status == 2'h2 | status == 2'h1; // @[BFS.scala 544:50]
  wire [31:0] _num_T_2 = num - 32'h4; // @[BFS.scala 560:18]
  wire [31:0] _num_T_6 = num > 32'h4 ? _num_T_2 : 32'h0; // @[BFS.scala 566:17]
  wire [31:0] _GEN_6 = r_demux_out_0_bits_rlast ? 32'h0 : _num_T_6; // @[BFS.scala 563:45 BFS.scala 564:11 BFS.scala 566:11]
  wire  _keep_0_T_3 = _T & r_demux_out_0_bits_rid[5]; // @[BFS.scala 573:33]
  wire  _keep_0_T_4 = num_regfile_io_dataOut > 32'h0; // @[BFS.scala 573:109]
  wire  _keep_0_T_6 = num > 32'h0; // @[BFS.scala 574:51]
  wire  _keep_0_T_10 = ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 575:36]
  wire  _keep_0_T_11 = _T & ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 575:33]
  wire [31:0] _keep_0_T_15 = r_demux_out_0_bits_rdata[63:32] + 32'h2; // @[BFS.scala 576:80]
  wire [2:0] _keep_0_T_22 = 3'h4 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_32 = {{29'd0}, _keep_0_T_22}; // @[BFS.scala 577:56]
  wire  _keep_0_T_23 = num > _GEN_32; // @[BFS.scala 577:56]
  wire  _keep_0_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_0_T_23; // @[Mux.scala 98:16]
  wire  _keep_0_T_26 = _T_8 ? _keep_0_T_6 : _keep_0_T_25; // @[Mux.scala 98:16]
  wire  keep_0 = _keep_0_T_3 ? _keep_0_T_4 : _keep_0_T_26; // @[Mux.scala 98:16]
  wire  _keep_1_T_4 = num_regfile_io_dataOut > 32'h1; // @[BFS.scala 573:109]
  wire  _keep_1_T_6 = num > 32'h1; // @[BFS.scala 574:51]
  wire [2:0] _keep_1_T_22 = 3'h5 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_33 = {{29'd0}, _keep_1_T_22}; // @[BFS.scala 577:56]
  wire  _keep_1_T_23 = num > _GEN_33; // @[BFS.scala 577:56]
  wire  _keep_1_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_1_T_23; // @[Mux.scala 98:16]
  wire  _keep_1_T_26 = _T_8 ? _keep_1_T_6 : _keep_1_T_25; // @[Mux.scala 98:16]
  wire  keep_1 = _keep_0_T_3 ? _keep_1_T_4 : _keep_1_T_26; // @[Mux.scala 98:16]
  wire  _keep_2_T_4 = num_regfile_io_dataOut > 32'h2; // @[BFS.scala 573:109]
  wire  _keep_2_T_6 = num > 32'h2; // @[BFS.scala 574:51]
  wire  _keep_2_T_16 = _keep_0_T_15 > 32'h2; // @[BFS.scala 576:87]
  wire [2:0] _keep_2_T_22 = 3'h6 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_34 = {{29'd0}, _keep_2_T_22}; // @[BFS.scala 577:56]
  wire  _keep_2_T_23 = num > _GEN_34; // @[BFS.scala 577:56]
  wire  _keep_2_T_25 = _keep_0_T_11 ? _keep_2_T_16 : _T_9 & _keep_2_T_23; // @[Mux.scala 98:16]
  wire  _keep_2_T_26 = _T_8 ? _keep_2_T_6 : _keep_2_T_25; // @[Mux.scala 98:16]
  wire  keep_2 = _keep_0_T_3 ? _keep_2_T_4 : _keep_2_T_26; // @[Mux.scala 98:16]
  wire  _keep_3_T_4 = num_regfile_io_dataOut > 32'h3; // @[BFS.scala 573:109]
  wire  _keep_3_T_6 = num > 32'h3; // @[BFS.scala 574:51]
  wire  _keep_3_T_16 = _keep_0_T_15 > 32'h3; // @[BFS.scala 576:87]
  wire [2:0] _keep_3_T_22 = 3'h7 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_35 = {{29'd0}, _keep_3_T_22}; // @[BFS.scala 577:56]
  wire  _keep_3_T_23 = num > _GEN_35; // @[BFS.scala 577:56]
  wire  _keep_3_T_25 = _keep_0_T_11 ? _keep_3_T_16 : _T_9 & _keep_3_T_23; // @[Mux.scala 98:16]
  wire  _keep_3_T_26 = _T_8 ? _keep_3_T_6 : _keep_3_T_25; // @[Mux.scala 98:16]
  wire  keep_3 = _keep_0_T_3 ? _keep_3_T_4 : _keep_3_T_26; // @[Mux.scala 98:16]
  wire [131:0] _vertex_out_fifo_io_din_T = {r_demux_out_0_bits_rdata,keep_3,keep_2,keep_1,keep_0}; // @[Cat.scala 30:58]
  reg  syncRecv_0; // @[BFS.scala 597:25]
  reg  syncRecv_1; // @[BFS.scala 597:25]
  reg  syncRecv_2; // @[BFS.scala 597:25]
  reg  syncRecv_3; // @[BFS.scala 597:25]
  reg  syncRecv_4; // @[BFS.scala 597:25]
  wire  _GEN_10 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_12 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_14 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_16 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_18 = io_recv_sync[4] | syncRecv_4; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 607:34]
  wire [31:0] _T_47 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_51 = _T_47[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_61 = vertex_out_fifo_data_count == 6'h0; // @[util.scala 211:19]
  wire  _T_62 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_61; // @[BFS.scala 612:71]
  wire [2:0] _GEN_21 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 621:53 BFS.scala 622:19 BFS.scala 466:30]
  wire [2:0] _GEN_22 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3 & syncRecv_4) ? 3'h0 :
    _GEN_21; // @[BFS.scala 615:71]
  wire  _T_79 = r_demux_out_0_valid & r_demux_out_0_ready & _keep_0_T_10; // @[BFS.scala 627:77]
  wire [63:0] _GEN_37 = {{32'd0}, r_demux_out_0_bits_rdata[63:32]}; // @[BFS.scala 629:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_37; // @[BFS.scala 629:46]
  wire  _T_82 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 632:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 636:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 638:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 472:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 481:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_free_ptr(edge_cache_io_free_ptr),
    .io_read_edge_num(edge_cache_io_read_edge_num),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_inflight_vtxs(edge_cache_io_inflight_vtxs)
  );
  r_demux r_demux ( // @[BFS.scala 485:23]
    .aclk(r_demux_aclk),
    .aresetn(r_demux_aresetn),
    .s_axis_tdata(r_demux_s_axis_tdata),
    .s_axis_tkeep(r_demux_s_axis_tkeep),
    .s_axis_tlast(r_demux_s_axis_tlast),
    .s_axis_tvalid(r_demux_s_axis_tvalid),
    .s_axis_tready(r_demux_s_axis_tready),
    .s_axis_tid(r_demux_s_axis_tid),
    .m_axis_tdata(r_demux_m_axis_tdata),
    .m_axis_tkeep(r_demux_m_axis_tkeep),
    .m_axis_tlast(r_demux_m_axis_tlast),
    .m_axis_tvalid(r_demux_m_axis_tvalid),
    .m_axis_tready(r_demux_m_axis_tready),
    .m_axis_tid(r_demux_m_axis_tid)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 506:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  regFile num_regfile ( // @[BFS.scala 519:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr),
    .io_wcount(num_regfile_io_wcount)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 581:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 507:13]
  assign io_ddr_r_ready = r_demux_s_axis_tready; // @[BFS.scala 494:18]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 477:52]
  assign io_xbar_out_valid = vertex_out_fifo_valid; // @[BFS.scala 584:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_dout[131:4]; // @[BFS.scala 586:52]
  assign io_xbar_out_bits_tkeep = vertex_out_fifo_dout[3:0]; // @[BFS.scala 585:52]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 469:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 607:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 476:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 475:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 515:80]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 473:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 474:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = r_demux_m_axis_tvalid[1]; // @[BFS.scala 497:42]
  assign edge_cache_io_in_bits_rdata = r_demux_m_axis_tdata[255:128]; // @[BFS.scala 500:46]
  assign edge_cache_io_in_bits_rid = r_demux_m_axis_tid[11:6]; // @[BFS.scala 498:42]
  assign edge_cache_io_in_bits_rlast = r_demux_m_axis_tlast[1]; // @[BFS.scala 499:46]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 516:17]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 483:32]
  assign edge_cache_io_free_ptr = num_regfile_io_wcount; // @[BFS.scala 524:26]
  assign edge_cache_io_inflight_vtxs = inflight_vtxs; // @[BFS.scala 484:31]
  assign r_demux_aclk = clock; // @[BFS.scala 492:34]
  assign r_demux_aresetn = ~reset; // @[BFS.scala 493:25]
  assign r_demux_s_axis_tdata = io_ddr_r_bits_rdata; // @[BFS.scala 488:27]
  assign r_demux_s_axis_tkeep = 16'hffff; // @[nf_arm_doce_top.scala 128:85]
  assign r_demux_s_axis_tlast = io_ddr_r_bits_rlast; // @[BFS.scala 489:27]
  assign r_demux_s_axis_tvalid = io_ddr_r_valid; // @[BFS.scala 487:28]
  assign r_demux_s_axis_tid = io_ddr_r_bits_rid; // @[BFS.scala 491:25]
  assign r_demux_m_axis_tready = {r_demux_out_1_ready,r_demux_out_0_ready}; // @[BFS.scala 503:84]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 516:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & inflight_vtxs < 64'h20; // @[BFS.scala 509:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_31; // @[BFS.scala 508:56]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id_lo}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 507:13]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = edge_cache_io_read_edge_num; // @[BFS.scala 522:25]
  assign num_regfile_io_writeFlag = arbi_io_in_0_ready & arbi_io_in_0_valid; // @[BFS.scala 520:51]
  assign num_regfile_io_rptr = r_demux_out_0_bits_rid[4:0]; // @[BFS.scala 369:7]
  assign num_regfile_io_wptr = num_regfile_io_wcount; // @[BFS.scala 521:23]
  assign vertex_out_fifo_din = _vertex_read_buffer_io_rd_en_T_2 ? 132'h800000001 : _vertex_out_fifo_io_din_T; // @[Mux.scala 98:16]
  assign vertex_out_fifo_wr_en = r_demux_out_0_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 589:52]
  assign vertex_out_fifo_rd_en = io_xbar_out_ready; // @[BFS.scala 588:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 583:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 582:42]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 466:30]
      upward_status <= 3'h0; // @[BFS.scala 466:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 608:57]
      upward_status <= 3'h1; // @[BFS.scala 609:19]
    end else if (upward_status == 3'h1 & (_T_51 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3 | syncRecv_4))
      ) begin // @[BFS.scala 610:105]
      upward_status <= 3'h2; // @[BFS.scala 611:19]
    end else if (_T_62 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 613:62]
      upward_status <= 3'h4; // @[BFS.scala 614:19]
    end else begin
      upward_status <= _GEN_22;
    end
    if (reset) begin // @[BFS.scala 467:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 467:30]
    end else if (!(_T_82 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 633:91]
      if (_T_82) begin // @[BFS.scala 635:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 636:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 637:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 638:19]
      end
    end
    if (reset) begin // @[BFS.scala 468:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 468:35]
    end else if (io_signal) begin // @[BFS.scala 625:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 626:24]
    end else if (_T_79 & _T) begin // @[BFS.scala 628:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 629:24]
    end
    if (reset) begin // @[BFS.scala 534:23]
      status <= 2'h0; // @[BFS.scala 534:23]
    end else if (status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 536:99]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 537:45]
        status <= 2'h0; // @[BFS.scala 538:14]
      end else if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 539:61]
        status <= 2'h2; // @[BFS.scala 540:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 542:14]
      end
    end else if (_T_10 & r_demux_out_0_valid & r_demux_out_0_ready & r_demux_out_0_bits_rlast) begin // @[BFS.scala 545:117]
      status <= 2'h0; // @[BFS.scala 546:14]
    end
    if (reset) begin // @[BFS.scala 535:20]
      num <= 32'h0; // @[BFS.scala 535:20]
    end else if (_T_4 & ~r_demux_out_0_bits_rlast) begin // @[BFS.scala 550:112]
      if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 551:55]
        num <= num_regfile_io_dataOut; // @[BFS.scala 552:11]
      end else begin
        num <= r_demux_out_0_bits_rdata[63:32]; // @[BFS.scala 554:11]
      end
    end else if (_T_8 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 556:114]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 557:45]
        num <= 32'h0; // @[BFS.scala 558:11]
      end else begin
        num <= _num_T_2; // @[BFS.scala 560:11]
      end
    end else if (_T_9 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 562:119]
      num <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_0 <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_1 <= _GEN_12;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_2 <= _GEN_14;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_3 <= _GEN_16;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_4 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_4 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_4 <= _GEN_18;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  status = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  num = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  syncRecv_4 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Broadcast_3(
  input          clock,
  input          reset,
  input          io_ddr_ar_ready,
  output         io_ddr_ar_valid,
  output [63:0]  io_ddr_ar_bits_araddr,
  output [5:0]   io_ddr_ar_bits_arid,
  output [7:0]   io_ddr_ar_bits_arlen,
  output [2:0]   io_ddr_ar_bits_arsize,
  output         io_ddr_r_ready,
  input          io_ddr_r_valid,
  input  [127:0] io_ddr_r_bits_rdata,
  input  [5:0]   io_ddr_r_bits_rid,
  input          io_ddr_r_bits_rlast,
  output         io_gather_in_ready,
  input          io_gather_in_valid,
  input  [31:0]  io_gather_in_bits_tdata,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [127:0] io_xbar_out_bits_tdata,
  output [3:0]   io_xbar_out_bits_tkeep,
  input  [63:0]  io_embedding_base_addr,
  input  [63:0]  io_edge_base_addr,
  input          io_signal,
  output [63:0]  io_traveled_edges,
  output         io_issue_sync,
  input  [4:0]   io_recv_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_read_buffer_full; // @[BFS.scala 472:34]
  wire [31:0] vertex_read_buffer_din; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_wr_en; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_empty; // @[BFS.scala 472:34]
  wire [31:0] vertex_read_buffer_dout; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_rd_en; // @[BFS.scala 472:34]
  wire [5:0] vertex_read_buffer_data_count; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_clk; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_srst; // @[BFS.scala 472:34]
  wire  vertex_read_buffer_valid; // @[BFS.scala 472:34]
  wire  edge_cache_clock; // @[BFS.scala 481:26]
  wire  edge_cache_reset; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_ready; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_valid; // @[BFS.scala 481:26]
  wire [127:0] edge_cache_io_in_bits_rdata; // @[BFS.scala 481:26]
  wire [5:0] edge_cache_io_in_bits_rid; // @[BFS.scala 481:26]
  wire  edge_cache_io_in_bits_rlast; // @[BFS.scala 481:26]
  wire  edge_cache_io_out_ready; // @[BFS.scala 481:26]
  wire  edge_cache_io_out_valid; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_out_bits_araddr; // @[BFS.scala 481:26]
  wire [5:0] edge_cache_io_out_bits_arid; // @[BFS.scala 481:26]
  wire [7:0] edge_cache_io_out_bits_arlen; // @[BFS.scala 481:26]
  wire [2:0] edge_cache_io_out_bits_arsize; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_edge_base_addr; // @[BFS.scala 481:26]
  wire [4:0] edge_cache_io_free_ptr; // @[BFS.scala 481:26]
  wire [31:0] edge_cache_io_read_edge_num; // @[BFS.scala 481:26]
  wire  edge_cache_io_read_edge_fifo_empty; // @[BFS.scala 481:26]
  wire [63:0] edge_cache_io_inflight_vtxs; // @[BFS.scala 481:26]
  wire  r_demux_aclk; // @[BFS.scala 485:23]
  wire  r_demux_aresetn; // @[BFS.scala 485:23]
  wire [127:0] r_demux_s_axis_tdata; // @[BFS.scala 485:23]
  wire [15:0] r_demux_s_axis_tkeep; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tlast; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tvalid; // @[BFS.scala 485:23]
  wire  r_demux_s_axis_tready; // @[BFS.scala 485:23]
  wire [5:0] r_demux_s_axis_tid; // @[BFS.scala 485:23]
  wire [255:0] r_demux_m_axis_tdata; // @[BFS.scala 485:23]
  wire [31:0] r_demux_m_axis_tkeep; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tlast; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tvalid; // @[BFS.scala 485:23]
  wire [1:0] r_demux_m_axis_tready; // @[BFS.scala 485:23]
  wire [11:0] r_demux_m_axis_tid; // @[BFS.scala 485:23]
  wire  arbi_clock; // @[BFS.scala 506:20]
  wire  arbi_reset; // @[BFS.scala 506:20]
  wire  arbi_io_in_0_ready; // @[BFS.scala 506:20]
  wire  arbi_io_in_0_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_in_0_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_in_0_bits_arid; // @[BFS.scala 506:20]
  wire [7:0] arbi_io_in_0_bits_arlen; // @[BFS.scala 506:20]
  wire [2:0] arbi_io_in_0_bits_arsize; // @[BFS.scala 506:20]
  wire  arbi_io_in_1_ready; // @[BFS.scala 506:20]
  wire  arbi_io_in_1_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_in_1_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_in_1_bits_arid; // @[BFS.scala 506:20]
  wire  arbi_io_out_ready; // @[BFS.scala 506:20]
  wire  arbi_io_out_valid; // @[BFS.scala 506:20]
  wire [63:0] arbi_io_out_bits_araddr; // @[BFS.scala 506:20]
  wire [5:0] arbi_io_out_bits_arid; // @[BFS.scala 506:20]
  wire [7:0] arbi_io_out_bits_arlen; // @[BFS.scala 506:20]
  wire [2:0] arbi_io_out_bits_arsize; // @[BFS.scala 506:20]
  wire  num_regfile_clock; // @[BFS.scala 519:27]
  wire  num_regfile_reset; // @[BFS.scala 519:27]
  wire [31:0] num_regfile_io_dataIn; // @[BFS.scala 519:27]
  wire [31:0] num_regfile_io_dataOut; // @[BFS.scala 519:27]
  wire  num_regfile_io_writeFlag; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_rptr; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_wptr; // @[BFS.scala 519:27]
  wire [4:0] num_regfile_io_wcount; // @[BFS.scala 519:27]
  wire  vertex_out_fifo_full; // @[BFS.scala 581:31]
  wire [131:0] vertex_out_fifo_din; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_wr_en; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_empty; // @[BFS.scala 581:31]
  wire [131:0] vertex_out_fifo_dout; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_rd_en; // @[BFS.scala 581:31]
  wire [5:0] vertex_out_fifo_data_count; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_clk; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_srst; // @[BFS.scala 581:31]
  wire  vertex_out_fifo_valid; // @[BFS.scala 581:31]
  (*dont_touch = "true" *)reg [2:0] upward_status; // @[BFS.scala 466:30]
  reg [63:0] inflight_vtxs; // @[BFS.scala 467:30]
  reg [63:0] traveled_edges_reg; // @[BFS.scala 468:35]
  wire [4:0] vertex_read_id_lo = vertex_read_buffer_data_count[4:0]; // @[BFS.scala 479:76 BFS.scala 479:76]
  wire  r_demux_out_0_valid = r_demux_m_axis_tvalid[0]; // @[BFS.scala 497:42]
  wire [5:0] r_demux_out_0_bits_rid = r_demux_m_axis_tid[5:0]; // @[BFS.scala 498:42]
  wire  r_demux_out_0_bits_rlast = r_demux_m_axis_tlast[0]; // @[BFS.scala 499:46]
  wire [127:0] r_demux_out_0_bits_rdata = r_demux_m_axis_tdata[127:0]; // @[BFS.scala 500:46]
  wire  r_demux_out_1_ready = edge_cache_io_in_ready; // @[BFS.scala 486:25 BFS.scala 504:20]
  wire  r_demux_out_0_ready = ~vertex_out_fifo_full; // @[BFS.scala 594:51]
  wire [37:0] _arbi_io_in_1_bits_araddr_T = {vertex_read_buffer_dout, 6'h0}; // @[BFS.scala 508:86]
  wire [63:0] _GEN_31 = {{26'd0}, _arbi_io_in_1_bits_araddr_T}; // @[BFS.scala 508:56]
  wire  _arbi_io_in_1_valid_T_3 = inflight_vtxs < 64'h20; // @[BFS.scala 509:116]
  wire  _vertex_read_buffer_io_rd_en_T_2 = upward_status == 3'h3; // @[BFS.scala 515:96]
  reg [1:0] status; // @[BFS.scala 534:23]
  reg [31:0] num; // @[BFS.scala 535:20]
  wire  _T = status == 2'h0; // @[BFS.scala 536:15]
  wire  _T_4 = status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready; // @[BFS.scala 536:66]
  wire  _T_8 = status == 2'h2; // @[BFS.scala 544:22]
  wire  _T_9 = status == 2'h1; // @[BFS.scala 544:60]
  wire  _T_10 = status == 2'h2 | status == 2'h1; // @[BFS.scala 544:50]
  wire [31:0] _num_T_2 = num - 32'h4; // @[BFS.scala 560:18]
  wire [31:0] _num_T_6 = num > 32'h4 ? _num_T_2 : 32'h0; // @[BFS.scala 566:17]
  wire [31:0] _GEN_6 = r_demux_out_0_bits_rlast ? 32'h0 : _num_T_6; // @[BFS.scala 563:45 BFS.scala 564:11 BFS.scala 566:11]
  wire  _keep_0_T_3 = _T & r_demux_out_0_bits_rid[5]; // @[BFS.scala 573:33]
  wire  _keep_0_T_4 = num_regfile_io_dataOut > 32'h0; // @[BFS.scala 573:109]
  wire  _keep_0_T_6 = num > 32'h0; // @[BFS.scala 574:51]
  wire  _keep_0_T_10 = ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 575:36]
  wire  _keep_0_T_11 = _T & ~r_demux_out_0_bits_rid[5]; // @[BFS.scala 575:33]
  wire [31:0] _keep_0_T_15 = r_demux_out_0_bits_rdata[63:32] + 32'h2; // @[BFS.scala 576:80]
  wire [2:0] _keep_0_T_22 = 3'h4 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_32 = {{29'd0}, _keep_0_T_22}; // @[BFS.scala 577:56]
  wire  _keep_0_T_23 = num > _GEN_32; // @[BFS.scala 577:56]
  wire  _keep_0_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_0_T_23; // @[Mux.scala 98:16]
  wire  _keep_0_T_26 = _T_8 ? _keep_0_T_6 : _keep_0_T_25; // @[Mux.scala 98:16]
  wire  keep_0 = _keep_0_T_3 ? _keep_0_T_4 : _keep_0_T_26; // @[Mux.scala 98:16]
  wire  _keep_1_T_4 = num_regfile_io_dataOut > 32'h1; // @[BFS.scala 573:109]
  wire  _keep_1_T_6 = num > 32'h1; // @[BFS.scala 574:51]
  wire [2:0] _keep_1_T_22 = 3'h5 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_33 = {{29'd0}, _keep_1_T_22}; // @[BFS.scala 577:56]
  wire  _keep_1_T_23 = num > _GEN_33; // @[BFS.scala 577:56]
  wire  _keep_1_T_25 = _keep_0_T_11 ? 1'h0 : _T_9 & _keep_1_T_23; // @[Mux.scala 98:16]
  wire  _keep_1_T_26 = _T_8 ? _keep_1_T_6 : _keep_1_T_25; // @[Mux.scala 98:16]
  wire  keep_1 = _keep_0_T_3 ? _keep_1_T_4 : _keep_1_T_26; // @[Mux.scala 98:16]
  wire  _keep_2_T_4 = num_regfile_io_dataOut > 32'h2; // @[BFS.scala 573:109]
  wire  _keep_2_T_6 = num > 32'h2; // @[BFS.scala 574:51]
  wire  _keep_2_T_16 = _keep_0_T_15 > 32'h2; // @[BFS.scala 576:87]
  wire [2:0] _keep_2_T_22 = 3'h6 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_34 = {{29'd0}, _keep_2_T_22}; // @[BFS.scala 577:56]
  wire  _keep_2_T_23 = num > _GEN_34; // @[BFS.scala 577:56]
  wire  _keep_2_T_25 = _keep_0_T_11 ? _keep_2_T_16 : _T_9 & _keep_2_T_23; // @[Mux.scala 98:16]
  wire  _keep_2_T_26 = _T_8 ? _keep_2_T_6 : _keep_2_T_25; // @[Mux.scala 98:16]
  wire  keep_2 = _keep_0_T_3 ? _keep_2_T_4 : _keep_2_T_26; // @[Mux.scala 98:16]
  wire  _keep_3_T_4 = num_regfile_io_dataOut > 32'h3; // @[BFS.scala 573:109]
  wire  _keep_3_T_6 = num > 32'h3; // @[BFS.scala 574:51]
  wire  _keep_3_T_16 = _keep_0_T_15 > 32'h3; // @[BFS.scala 576:87]
  wire [2:0] _keep_3_T_22 = 3'h7 - 3'h2; // @[BFS.scala 577:78]
  wire [31:0] _GEN_35 = {{29'd0}, _keep_3_T_22}; // @[BFS.scala 577:56]
  wire  _keep_3_T_23 = num > _GEN_35; // @[BFS.scala 577:56]
  wire  _keep_3_T_25 = _keep_0_T_11 ? _keep_3_T_16 : _T_9 & _keep_3_T_23; // @[Mux.scala 98:16]
  wire  _keep_3_T_26 = _T_8 ? _keep_3_T_6 : _keep_3_T_25; // @[Mux.scala 98:16]
  wire  keep_3 = _keep_0_T_3 ? _keep_3_T_4 : _keep_3_T_26; // @[Mux.scala 98:16]
  wire [131:0] _vertex_out_fifo_io_din_T = {r_demux_out_0_bits_rdata,keep_3,keep_2,keep_1,keep_0}; // @[Cat.scala 30:58]
  reg  syncRecv_0; // @[BFS.scala 597:25]
  reg  syncRecv_1; // @[BFS.scala 597:25]
  reg  syncRecv_2; // @[BFS.scala 597:25]
  reg  syncRecv_3; // @[BFS.scala 597:25]
  reg  syncRecv_4; // @[BFS.scala 597:25]
  wire  _GEN_10 = io_recv_sync[0] | syncRecv_0; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_12 = io_recv_sync[1] | syncRecv_1; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_14 = io_recv_sync[2] | syncRecv_2; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_16 = io_recv_sync[3] | syncRecv_3; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _GEN_18 = io_recv_sync[4] | syncRecv_4; // @[BFS.scala 602:34 BFS.scala 603:11 BFS.scala 597:25]
  wire  _io_issue_sync_T = upward_status == 3'h4; // @[BFS.scala 607:34]
  wire [31:0] _T_47 = {{31'd0}, vertex_read_buffer_dout[31]}; // @[util.scala 207:12]
  wire  _T_51 = _T_47[0] & ~vertex_read_buffer_empty; // @[util.scala 207:36]
  wire  _T_61 = vertex_out_fifo_data_count == 6'h0; // @[util.scala 211:19]
  wire  _T_62 = upward_status == 3'h2 & inflight_vtxs == 64'h0 & _T_61; // @[BFS.scala 612:71]
  wire [2:0] _GEN_21 = _vertex_read_buffer_io_rd_en_T_2 ? 3'h0 : upward_status; // @[BFS.scala 621:53 BFS.scala 622:19 BFS.scala 466:30]
  wire [2:0] _GEN_22 = _io_issue_sync_T & (syncRecv_0 & syncRecv_1 & syncRecv_2 & syncRecv_3 & syncRecv_4) ? 3'h0 :
    _GEN_21; // @[BFS.scala 615:71]
  wire  _T_79 = r_demux_out_0_valid & r_demux_out_0_ready & _keep_0_T_10; // @[BFS.scala 627:77]
  wire [63:0] _GEN_37 = {{32'd0}, r_demux_out_0_bits_rdata[63:32]}; // @[BFS.scala 629:46]
  wire [63:0] _traveled_edges_reg_T_2 = traveled_edges_reg + _GEN_37; // @[BFS.scala 629:46]
  wire  _T_82 = io_ddr_ar_valid & io_ddr_ar_ready; // @[BFS.scala 632:24]
  wire [63:0] _inflight_vtxs_T_1 = inflight_vtxs + 64'h1; // @[BFS.scala 636:36]
  wire [63:0] _inflight_vtxs_T_3 = inflight_vtxs - 64'h1; // @[BFS.scala 638:36]
  vid_fifo vertex_read_buffer ( // @[BFS.scala 472:34]
    .full(vertex_read_buffer_full),
    .din(vertex_read_buffer_din),
    .wr_en(vertex_read_buffer_wr_en),
    .empty(vertex_read_buffer_empty),
    .dout(vertex_read_buffer_dout),
    .rd_en(vertex_read_buffer_rd_en),
    .data_count(vertex_read_buffer_data_count),
    .clk(vertex_read_buffer_clk),
    .srst(vertex_read_buffer_srst),
    .valid(vertex_read_buffer_valid)
  );
  readEdge_engine edge_cache ( // @[BFS.scala 481:26]
    .clock(edge_cache_clock),
    .reset(edge_cache_reset),
    .io_in_ready(edge_cache_io_in_ready),
    .io_in_valid(edge_cache_io_in_valid),
    .io_in_bits_rdata(edge_cache_io_in_bits_rdata),
    .io_in_bits_rid(edge_cache_io_in_bits_rid),
    .io_in_bits_rlast(edge_cache_io_in_bits_rlast),
    .io_out_ready(edge_cache_io_out_ready),
    .io_out_valid(edge_cache_io_out_valid),
    .io_out_bits_araddr(edge_cache_io_out_bits_araddr),
    .io_out_bits_arid(edge_cache_io_out_bits_arid),
    .io_out_bits_arlen(edge_cache_io_out_bits_arlen),
    .io_out_bits_arsize(edge_cache_io_out_bits_arsize),
    .io_edge_base_addr(edge_cache_io_edge_base_addr),
    .io_free_ptr(edge_cache_io_free_ptr),
    .io_read_edge_num(edge_cache_io_read_edge_num),
    .io_read_edge_fifo_empty(edge_cache_io_read_edge_fifo_empty),
    .io_inflight_vtxs(edge_cache_io_inflight_vtxs)
  );
  r_demux r_demux ( // @[BFS.scala 485:23]
    .aclk(r_demux_aclk),
    .aresetn(r_demux_aresetn),
    .s_axis_tdata(r_demux_s_axis_tdata),
    .s_axis_tkeep(r_demux_s_axis_tkeep),
    .s_axis_tlast(r_demux_s_axis_tlast),
    .s_axis_tvalid(r_demux_s_axis_tvalid),
    .s_axis_tready(r_demux_s_axis_tready),
    .s_axis_tid(r_demux_s_axis_tid),
    .m_axis_tdata(r_demux_m_axis_tdata),
    .m_axis_tkeep(r_demux_m_axis_tkeep),
    .m_axis_tlast(r_demux_m_axis_tlast),
    .m_axis_tvalid(r_demux_m_axis_tvalid),
    .m_axis_tready(r_demux_m_axis_tready),
    .m_axis_tid(r_demux_m_axis_tid)
  );
  AMBA_Arbiter arbi ( // @[BFS.scala 506:20]
    .clock(arbi_clock),
    .reset(arbi_reset),
    .io_in_0_ready(arbi_io_in_0_ready),
    .io_in_0_valid(arbi_io_in_0_valid),
    .io_in_0_bits_araddr(arbi_io_in_0_bits_araddr),
    .io_in_0_bits_arid(arbi_io_in_0_bits_arid),
    .io_in_0_bits_arlen(arbi_io_in_0_bits_arlen),
    .io_in_0_bits_arsize(arbi_io_in_0_bits_arsize),
    .io_in_1_ready(arbi_io_in_1_ready),
    .io_in_1_valid(arbi_io_in_1_valid),
    .io_in_1_bits_araddr(arbi_io_in_1_bits_araddr),
    .io_in_1_bits_arid(arbi_io_in_1_bits_arid),
    .io_out_ready(arbi_io_out_ready),
    .io_out_valid(arbi_io_out_valid),
    .io_out_bits_araddr(arbi_io_out_bits_araddr),
    .io_out_bits_arid(arbi_io_out_bits_arid),
    .io_out_bits_arlen(arbi_io_out_bits_arlen),
    .io_out_bits_arsize(arbi_io_out_bits_arsize)
  );
  regFile num_regfile ( // @[BFS.scala 519:27]
    .clock(num_regfile_clock),
    .reset(num_regfile_reset),
    .io_dataIn(num_regfile_io_dataIn),
    .io_dataOut(num_regfile_io_dataOut),
    .io_writeFlag(num_regfile_io_writeFlag),
    .io_rptr(num_regfile_io_rptr),
    .io_wptr(num_regfile_io_wptr),
    .io_wcount(num_regfile_io_wcount)
  );
  edge_fifo vertex_out_fifo ( // @[BFS.scala 581:31]
    .full(vertex_out_fifo_full),
    .din(vertex_out_fifo_din),
    .wr_en(vertex_out_fifo_wr_en),
    .empty(vertex_out_fifo_empty),
    .dout(vertex_out_fifo_dout),
    .rd_en(vertex_out_fifo_rd_en),
    .data_count(vertex_out_fifo_data_count),
    .clk(vertex_out_fifo_clk),
    .srst(vertex_out_fifo_srst),
    .valid(vertex_out_fifo_valid)
  );
  assign io_ddr_ar_valid = arbi_io_out_valid; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_araddr = arbi_io_out_bits_araddr; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arid = arbi_io_out_bits_arid; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arlen = arbi_io_out_bits_arlen; // @[BFS.scala 507:13]
  assign io_ddr_ar_bits_arsize = arbi_io_out_bits_arsize; // @[BFS.scala 507:13]
  assign io_ddr_r_ready = r_demux_s_axis_tready; // @[BFS.scala 494:18]
  assign io_gather_in_ready = ~vertex_read_buffer_full; // @[BFS.scala 477:52]
  assign io_xbar_out_valid = vertex_out_fifo_valid; // @[BFS.scala 584:21]
  assign io_xbar_out_bits_tdata = vertex_out_fifo_dout[131:4]; // @[BFS.scala 586:52]
  assign io_xbar_out_bits_tkeep = vertex_out_fifo_dout[3:0]; // @[BFS.scala 585:52]
  assign io_traveled_edges = traveled_edges_reg; // @[BFS.scala 469:21]
  assign io_issue_sync = upward_status == 3'h4; // @[BFS.scala 607:34]
  assign vertex_read_buffer_din = io_gather_in_bits_tdata; // @[BFS.scala 476:29]
  assign vertex_read_buffer_wr_en = io_gather_in_valid; // @[BFS.scala 475:31]
  assign vertex_read_buffer_rd_en = arbi_io_in_1_ready & _arbi_io_in_1_valid_T_3 | upward_status == 3'h3; // @[BFS.scala 515:80]
  assign vertex_read_buffer_clk = clock; // @[BFS.scala 473:44]
  assign vertex_read_buffer_srst = reset; // @[BFS.scala 474:45]
  assign edge_cache_clock = clock;
  assign edge_cache_reset = reset;
  assign edge_cache_io_in_valid = r_demux_m_axis_tvalid[1]; // @[BFS.scala 497:42]
  assign edge_cache_io_in_bits_rdata = r_demux_m_axis_tdata[255:128]; // @[BFS.scala 500:46]
  assign edge_cache_io_in_bits_rid = r_demux_m_axis_tid[11:6]; // @[BFS.scala 498:42]
  assign edge_cache_io_in_bits_rlast = r_demux_m_axis_tlast[1]; // @[BFS.scala 499:46]
  assign edge_cache_io_out_ready = arbi_io_in_0_ready; // @[BFS.scala 516:17]
  assign edge_cache_io_edge_base_addr = io_edge_base_addr; // @[BFS.scala 483:32]
  assign edge_cache_io_free_ptr = num_regfile_io_wcount; // @[BFS.scala 524:26]
  assign edge_cache_io_inflight_vtxs = inflight_vtxs; // @[BFS.scala 484:31]
  assign r_demux_aclk = clock; // @[BFS.scala 492:34]
  assign r_demux_aresetn = ~reset; // @[BFS.scala 493:25]
  assign r_demux_s_axis_tdata = io_ddr_r_bits_rdata; // @[BFS.scala 488:27]
  assign r_demux_s_axis_tkeep = 16'hffff; // @[nf_arm_doce_top.scala 128:85]
  assign r_demux_s_axis_tlast = io_ddr_r_bits_rlast; // @[BFS.scala 489:27]
  assign r_demux_s_axis_tvalid = io_ddr_r_valid; // @[BFS.scala 487:28]
  assign r_demux_s_axis_tid = io_ddr_r_bits_rid; // @[BFS.scala 491:25]
  assign r_demux_m_axis_tready = {r_demux_out_1_ready,r_demux_out_0_ready}; // @[BFS.scala 503:84]
  assign arbi_clock = clock;
  assign arbi_reset = reset;
  assign arbi_io_in_0_valid = edge_cache_io_out_valid; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_araddr = edge_cache_io_out_bits_araddr; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arid = edge_cache_io_out_bits_arid; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arlen = edge_cache_io_out_bits_arlen; // @[BFS.scala 516:17]
  assign arbi_io_in_0_bits_arsize = edge_cache_io_out_bits_arsize; // @[BFS.scala 516:17]
  assign arbi_io_in_1_valid = vertex_read_buffer_valid & ~vertex_read_buffer_dout[31] & inflight_vtxs < 64'h20; // @[BFS.scala 509:99]
  assign arbi_io_in_1_bits_araddr = io_embedding_base_addr + _GEN_31; // @[BFS.scala 508:56]
  assign arbi_io_in_1_bits_arid = {1'h0,vertex_read_id_lo}; // @[Cat.scala 30:58]
  assign arbi_io_out_ready = io_ddr_ar_ready; // @[BFS.scala 507:13]
  assign num_regfile_clock = clock;
  assign num_regfile_reset = reset;
  assign num_regfile_io_dataIn = edge_cache_io_read_edge_num; // @[BFS.scala 522:25]
  assign num_regfile_io_writeFlag = arbi_io_in_0_ready & arbi_io_in_0_valid; // @[BFS.scala 520:51]
  assign num_regfile_io_rptr = r_demux_out_0_bits_rid[4:0]; // @[BFS.scala 369:7]
  assign num_regfile_io_wptr = num_regfile_io_wcount; // @[BFS.scala 521:23]
  assign vertex_out_fifo_din = _vertex_read_buffer_io_rd_en_T_2 ? 132'h800000001 : _vertex_out_fifo_io_din_T; // @[Mux.scala 98:16]
  assign vertex_out_fifo_wr_en = r_demux_out_0_valid | _vertex_read_buffer_io_rd_en_T_2; // @[BFS.scala 589:52]
  assign vertex_out_fifo_rd_en = io_xbar_out_ready; // @[BFS.scala 588:28]
  assign vertex_out_fifo_clk = clock; // @[BFS.scala 583:41]
  assign vertex_out_fifo_srst = reset; // @[BFS.scala 582:42]
  always @(posedge clock) begin
    if (reset) begin // @[BFS.scala 466:30]
      upward_status <= 3'h0; // @[BFS.scala 466:30]
    end else if (io_signal & upward_status == 3'h0) begin // @[BFS.scala 608:57]
      upward_status <= 3'h1; // @[BFS.scala 609:19]
    end else if (upward_status == 3'h1 & (_T_51 | (syncRecv_0 | syncRecv_1 | syncRecv_2 | syncRecv_3 | syncRecv_4))
      ) begin // @[BFS.scala 610:105]
      upward_status <= 3'h2; // @[BFS.scala 611:19]
    end else if (_T_62 & edge_cache_io_read_edge_fifo_empty) begin // @[BFS.scala 613:62]
      upward_status <= 3'h4; // @[BFS.scala 614:19]
    end else begin
      upward_status <= _GEN_22;
    end
    if (reset) begin // @[BFS.scala 467:30]
      inflight_vtxs <= 64'h0; // @[BFS.scala 467:30]
    end else if (!(_T_82 & io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast)) begin // @[BFS.scala 633:91]
      if (_T_82) begin // @[BFS.scala 635:49]
        inflight_vtxs <= _inflight_vtxs_T_1; // @[BFS.scala 636:19]
      end else if (io_ddr_r_valid & io_ddr_r_ready & io_ddr_r_bits_rlast) begin // @[BFS.scala 637:97]
        inflight_vtxs <= _inflight_vtxs_T_3; // @[BFS.scala 638:19]
      end
    end
    if (reset) begin // @[BFS.scala 468:35]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 468:35]
    end else if (io_signal) begin // @[BFS.scala 625:18]
      traveled_edges_reg <= 64'h0; // @[BFS.scala 626:24]
    end else if (_T_79 & _T) begin // @[BFS.scala 628:33]
      traveled_edges_reg <= _traveled_edges_reg_T_2; // @[BFS.scala 629:24]
    end
    if (reset) begin // @[BFS.scala 534:23]
      status <= 2'h0; // @[BFS.scala 534:23]
    end else if (status == 2'h0 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 536:99]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 537:45]
        status <= 2'h0; // @[BFS.scala 538:14]
      end else if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 539:61]
        status <= 2'h2; // @[BFS.scala 540:14]
      end else begin
        status <= 2'h1; // @[BFS.scala 542:14]
      end
    end else if (_T_10 & r_demux_out_0_valid & r_demux_out_0_ready & r_demux_out_0_bits_rlast) begin // @[BFS.scala 545:117]
      status <= 2'h0; // @[BFS.scala 546:14]
    end
    if (reset) begin // @[BFS.scala 535:20]
      num <= 32'h0; // @[BFS.scala 535:20]
    end else if (_T_4 & ~r_demux_out_0_bits_rlast) begin // @[BFS.scala 550:112]
      if (r_demux_out_0_bits_rid[5]) begin // @[BFS.scala 551:55]
        num <= num_regfile_io_dataOut; // @[BFS.scala 552:11]
      end else begin
        num <= r_demux_out_0_bits_rdata[63:32]; // @[BFS.scala 554:11]
      end
    end else if (_T_8 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 556:114]
      if (r_demux_out_0_bits_rlast) begin // @[BFS.scala 557:45]
        num <= 32'h0; // @[BFS.scala 558:11]
      end else begin
        num <= _num_T_2; // @[BFS.scala 560:11]
      end
    end else if (_T_9 & r_demux_out_0_valid & r_demux_out_0_ready) begin // @[BFS.scala 562:119]
      num <= _GEN_6;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_0 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_0 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_0 <= _GEN_10;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_1 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_1 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_1 <= _GEN_12;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_2 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_2 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_2 <= _GEN_14;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_3 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_3 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_3 <= _GEN_16;
    end
    if (reset) begin // @[BFS.scala 597:25]
      syncRecv_4 <= 1'h0; // @[BFS.scala 597:25]
    end else if (io_signal) begin // @[BFS.scala 600:22]
      syncRecv_4 <= 1'h0; // @[BFS.scala 601:11]
    end else begin
      syncRecv_4 <= _GEN_18;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  upward_status = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  inflight_vtxs = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  traveled_edges_reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  status = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  num = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  syncRecv_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  syncRecv_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  syncRecv_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  syncRecv_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  syncRecv_4 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Remote_xbar(
  input           clock,
  input           reset,
  output          io_ddr_in_0_ready,
  input           io_ddr_in_0_valid,
  input  [127:0]  io_ddr_in_0_bits_tdata,
  input  [3:0]    io_ddr_in_0_bits_tkeep,
  output          io_ddr_in_1_ready,
  input           io_ddr_in_1_valid,
  input  [127:0]  io_ddr_in_1_bits_tdata,
  input  [3:0]    io_ddr_in_1_bits_tkeep,
  output          io_ddr_in_2_ready,
  input           io_ddr_in_2_valid,
  input  [127:0]  io_ddr_in_2_bits_tdata,
  input  [3:0]    io_ddr_in_2_bits_tkeep,
  output          io_ddr_in_3_ready,
  input           io_ddr_in_3_valid,
  input  [127:0]  io_ddr_in_3_bits_tdata,
  input  [3:0]    io_ddr_in_3_bits_tkeep,
  input           io_pe_out_0_ready,
  output          io_pe_out_0_valid,
  output [1023:0] io_pe_out_0_bits_tdata,
  output [31:0]   io_pe_out_0_bits_tkeep,
  input           io_pe_out_1_ready,
  output          io_pe_out_1_valid,
  output [1023:0] io_pe_out_1_bits_tdata,
  output [31:0]   io_pe_out_1_bits_tkeep,
  input           io_pe_out_2_ready,
  output          io_pe_out_2_valid,
  output [1023:0] io_pe_out_2_bits_tdata,
  output [31:0]   io_pe_out_2_bits_tkeep,
  input           io_pe_out_3_ready,
  output          io_pe_out_3_valid,
  output [1023:0] io_pe_out_3_bits_tdata,
  output [31:0]   io_pe_out_3_bits_tkeep,
  input           io_pe_out_4_ready,
  output          io_pe_out_4_valid,
  output [1023:0] io_pe_out_4_bits_tdata,
  output [31:0]   io_pe_out_4_bits_tkeep,
  input           io_pe_out_5_ready,
  output          io_pe_out_5_valid,
  output [1023:0] io_pe_out_5_bits_tdata,
  output [31:0]   io_pe_out_5_bits_tkeep,
  input           io_pe_out_6_ready,
  output          io_pe_out_6_valid,
  output [1023:0] io_pe_out_6_bits_tdata,
  output [31:0]   io_pe_out_6_bits_tkeep,
  input           io_pe_out_7_ready,
  output          io_pe_out_7_valid,
  output [1023:0] io_pe_out_7_bits_tdata,
  output [31:0]   io_pe_out_7_bits_tkeep,
  input           io_pe_out_8_ready,
  output          io_pe_out_8_valid,
  output [1023:0] io_pe_out_8_bits_tdata,
  output [31:0]   io_pe_out_8_bits_tkeep,
  input           io_pe_out_9_ready,
  output          io_pe_out_9_valid,
  output [1023:0] io_pe_out_9_bits_tdata,
  output [31:0]   io_pe_out_9_bits_tkeep,
  input           io_pe_out_10_ready,
  output          io_pe_out_10_valid,
  output [1023:0] io_pe_out_10_bits_tdata,
  output [31:0]   io_pe_out_10_bits_tkeep,
  input           io_pe_out_11_ready,
  output          io_pe_out_11_valid,
  output [1023:0] io_pe_out_11_bits_tdata,
  output [31:0]   io_pe_out_11_bits_tkeep,
  input           io_pe_out_12_ready,
  output          io_pe_out_12_valid,
  output [1023:0] io_pe_out_12_bits_tdata,
  output [31:0]   io_pe_out_12_bits_tkeep,
  input           io_pe_out_13_ready,
  output          io_pe_out_13_valid,
  output [1023:0] io_pe_out_13_bits_tdata,
  output [31:0]   io_pe_out_13_bits_tkeep,
  input           io_pe_out_14_ready,
  output          io_pe_out_14_valid,
  output [1023:0] io_pe_out_14_bits_tdata,
  output [31:0]   io_pe_out_14_bits_tkeep,
  input           io_pe_out_15_ready,
  output          io_pe_out_15_valid,
  output [1023:0] io_pe_out_15_bits_tdata,
  output [31:0]   io_pe_out_15_bits_tkeep,
  input           io_remote_out_ready,
  output          io_remote_out_valid,
  output [511:0]  io_remote_out_bits_tdata,
  output [15:0]   io_remote_out_bits_tkeep,
  output          io_remote_in_ready,
  input           io_remote_in_valid,
  input  [511:0]  io_remote_in_bits_tdata,
  input  [15:0]   io_remote_in_bits_tkeep
);
  wire  combiner_level0_aclk; // @[bfs_remote.scala 238:31]
  wire  combiner_level0_aresetn; // @[bfs_remote.scala 238:31]
  wire [511:0] combiner_level0_s_axis_tdata; // @[bfs_remote.scala 238:31]
  wire [63:0] combiner_level0_s_axis_tkeep; // @[bfs_remote.scala 238:31]
  wire [3:0] combiner_level0_s_axis_tlast; // @[bfs_remote.scala 238:31]
  wire [3:0] combiner_level0_s_axis_tvalid; // @[bfs_remote.scala 238:31]
  wire [3:0] combiner_level0_s_axis_tready; // @[bfs_remote.scala 238:31]
  wire [3:0] combiner_level0_s_axis_tid; // @[bfs_remote.scala 238:31]
  wire [511:0] combiner_level0_m_axis_tdata; // @[bfs_remote.scala 238:31]
  wire [63:0] combiner_level0_m_axis_tkeep; // @[bfs_remote.scala 238:31]
  wire  combiner_level0_m_axis_tlast; // @[bfs_remote.scala 238:31]
  wire  combiner_level0_m_axis_tvalid; // @[bfs_remote.scala 238:31]
  wire  combiner_level0_m_axis_tready; // @[bfs_remote.scala 238:31]
  wire  combiner_level0_m_axis_tid; // @[bfs_remote.scala 238:31]
  wire  xbar_level0_aclk; // @[bfs_remote.scala 250:27]
  wire  xbar_level0_aresetn; // @[bfs_remote.scala 250:27]
  wire [511:0] xbar_level0_s_axis_tdata; // @[bfs_remote.scala 250:27]
  wire [63:0] xbar_level0_s_axis_tkeep; // @[bfs_remote.scala 250:27]
  wire  xbar_level0_s_axis_tlast; // @[bfs_remote.scala 250:27]
  wire  xbar_level0_s_axis_tvalid; // @[bfs_remote.scala 250:27]
  wire  xbar_level0_s_axis_tready; // @[bfs_remote.scala 250:27]
  wire  xbar_level0_s_axis_tid; // @[bfs_remote.scala 250:27]
  wire [1023:0] xbar_level0_m_axis_tdata; // @[bfs_remote.scala 250:27]
  wire [127:0] xbar_level0_m_axis_tkeep; // @[bfs_remote.scala 250:27]
  wire [1:0] xbar_level0_m_axis_tlast; // @[bfs_remote.scala 250:27]
  wire [1:0] xbar_level0_m_axis_tvalid; // @[bfs_remote.scala 250:27]
  wire [1:0] xbar_level0_m_axis_tready; // @[bfs_remote.scala 250:27]
  wire [1:0] xbar_level0_m_axis_tid; // @[bfs_remote.scala 250:27]
  wire  combiner_level1_aclk; // @[bfs_remote.scala 257:31]
  wire  combiner_level1_aresetn; // @[bfs_remote.scala 257:31]
  wire [1023:0] combiner_level1_s_axis_tdata; // @[bfs_remote.scala 257:31]
  wire [127:0] combiner_level1_s_axis_tkeep; // @[bfs_remote.scala 257:31]
  wire [1:0] combiner_level1_s_axis_tlast; // @[bfs_remote.scala 257:31]
  wire [1:0] combiner_level1_s_axis_tvalid; // @[bfs_remote.scala 257:31]
  wire [1:0] combiner_level1_s_axis_tready; // @[bfs_remote.scala 257:31]
  wire [1:0] combiner_level1_s_axis_tid; // @[bfs_remote.scala 257:31]
  wire [1023:0] combiner_level1_m_axis_tdata; // @[bfs_remote.scala 257:31]
  wire [127:0] combiner_level1_m_axis_tkeep; // @[bfs_remote.scala 257:31]
  wire  combiner_level1_m_axis_tlast; // @[bfs_remote.scala 257:31]
  wire  combiner_level1_m_axis_tvalid; // @[bfs_remote.scala 257:31]
  wire  combiner_level1_m_axis_tready; // @[bfs_remote.scala 257:31]
  wire  combiner_level1_m_axis_tid; // @[bfs_remote.scala 257:31]
  wire  xbar_level1_aclk; // @[bfs_remote.scala 268:27]
  wire  xbar_level1_aresetn; // @[bfs_remote.scala 268:27]
  wire [1023:0] xbar_level1_s_axis_tdata; // @[bfs_remote.scala 268:27]
  wire [127:0] xbar_level1_s_axis_tkeep; // @[bfs_remote.scala 268:27]
  wire  xbar_level1_s_axis_tlast; // @[bfs_remote.scala 268:27]
  wire  xbar_level1_s_axis_tvalid; // @[bfs_remote.scala 268:27]
  wire  xbar_level1_s_axis_tready; // @[bfs_remote.scala 268:27]
  wire  xbar_level1_s_axis_tid; // @[bfs_remote.scala 268:27]
  wire [16383:0] xbar_level1_m_axis_tdata; // @[bfs_remote.scala 268:27]
  wire [2047:0] xbar_level1_m_axis_tkeep; // @[bfs_remote.scala 268:27]
  wire [15:0] xbar_level1_m_axis_tlast; // @[bfs_remote.scala 268:27]
  wire [15:0] xbar_level1_m_axis_tvalid; // @[bfs_remote.scala 268:27]
  wire [15:0] xbar_level1_m_axis_tready; // @[bfs_remote.scala 268:27]
  wire [15:0] xbar_level1_m_axis_tid; // @[bfs_remote.scala 268:27]
  wire [255:0] combiner_level0_io_s_axis_tdata_lo = {io_ddr_in_1_bits_tdata,io_ddr_in_0_bits_tdata}; // @[bfs_remote.scala 241:103]
  wire [255:0] combiner_level0_io_s_axis_tdata_hi = {io_ddr_in_3_bits_tdata,io_ddr_in_2_bits_tdata}; // @[bfs_remote.scala 241:103]
  wire  _combiner_level0_io_s_axis_tkeep_T_4 = io_ddr_in_0_bits_tkeep[0] & io_ddr_in_0_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_5 = io_ddr_in_0_bits_tkeep[1] & io_ddr_in_0_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_6 = io_ddr_in_0_bits_tkeep[2] & io_ddr_in_0_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_7 = io_ddr_in_0_bits_tkeep[3] & io_ddr_in_0_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_12 = io_ddr_in_1_bits_tkeep[0] & io_ddr_in_1_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_13 = io_ddr_in_1_bits_tkeep[1] & io_ddr_in_1_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_14 = io_ddr_in_1_bits_tkeep[2] & io_ddr_in_1_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_15 = io_ddr_in_1_bits_tkeep[3] & io_ddr_in_1_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_20 = io_ddr_in_2_bits_tkeep[0] & io_ddr_in_2_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_21 = io_ddr_in_2_bits_tkeep[1] & io_ddr_in_2_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_22 = io_ddr_in_2_bits_tkeep[2] & io_ddr_in_2_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_23 = io_ddr_in_2_bits_tkeep[3] & io_ddr_in_2_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_28 = io_ddr_in_3_bits_tkeep[0] & io_ddr_in_3_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_29 = io_ddr_in_3_bits_tkeep[1] & io_ddr_in_3_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_30 = io_ddr_in_3_bits_tkeep[2] & io_ddr_in_3_valid; // @[bfs_remote.scala 242:125]
  wire  _combiner_level0_io_s_axis_tkeep_T_31 = io_ddr_in_3_bits_tkeep[3] & io_ddr_in_3_valid; // @[bfs_remote.scala 242:125]
  wire [7:0] combiner_level0_io_s_axis_tkeep_lo = {_combiner_level0_io_s_axis_tkeep_T_15,
    _combiner_level0_io_s_axis_tkeep_T_14,_combiner_level0_io_s_axis_tkeep_T_13,_combiner_level0_io_s_axis_tkeep_T_12,
    _combiner_level0_io_s_axis_tkeep_T_7,_combiner_level0_io_s_axis_tkeep_T_6,_combiner_level0_io_s_axis_tkeep_T_5,
    _combiner_level0_io_s_axis_tkeep_T_4}; // @[bfs_remote.scala 243:33]
  wire [15:0] _combiner_level0_io_s_axis_tkeep_T_32 = {_combiner_level0_io_s_axis_tkeep_T_31,
    _combiner_level0_io_s_axis_tkeep_T_30,_combiner_level0_io_s_axis_tkeep_T_29,_combiner_level0_io_s_axis_tkeep_T_28,
    _combiner_level0_io_s_axis_tkeep_T_23,_combiner_level0_io_s_axis_tkeep_T_22,_combiner_level0_io_s_axis_tkeep_T_21,
    _combiner_level0_io_s_axis_tkeep_T_20,combiner_level0_io_s_axis_tkeep_lo}; // @[bfs_remote.scala 243:33]
  wire  _combiner_level0_io_s_axis_tvalid_T_2 = io_ddr_in_0_valid | io_ddr_in_1_valid | io_ddr_in_2_valid |
    io_ddr_in_3_valid; // @[bfs_remote.scala 245:104]
  wire [1:0] combiner_level0_io_s_axis_tvalid_lo = {_combiner_level0_io_s_axis_tvalid_T_2,
    _combiner_level0_io_s_axis_tvalid_T_2}; // @[bfs_remote.scala 245:116]
  wire [511:0] combiner_level1_io_s_axis_tdata_hi = xbar_level0_m_axis_tdata[511:0]; // @[bfs_remote.scala 260:69]
  wire [63:0] combiner_level1_io_s_axis_tkeep_hi = xbar_level0_m_axis_tkeep[63:0]; // @[bfs_remote.scala 261:69]
  wire  _combiner_level1_io_s_axis_tkeep_T_16 = io_remote_in_bits_tkeep[0] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_17 = io_remote_in_bits_tkeep[1] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_18 = io_remote_in_bits_tkeep[2] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_19 = io_remote_in_bits_tkeep[3] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_20 = io_remote_in_bits_tkeep[4] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_21 = io_remote_in_bits_tkeep[5] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_22 = io_remote_in_bits_tkeep[6] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_23 = io_remote_in_bits_tkeep[7] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_24 = io_remote_in_bits_tkeep[8] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_25 = io_remote_in_bits_tkeep[9] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_26 = io_remote_in_bits_tkeep[10] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_27 = io_remote_in_bits_tkeep[11] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_28 = io_remote_in_bits_tkeep[12] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_29 = io_remote_in_bits_tkeep[13] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_30 = io_remote_in_bits_tkeep[14] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire  _combiner_level1_io_s_axis_tkeep_T_31 = io_remote_in_bits_tkeep[15] & io_remote_in_valid; // @[bfs_remote.scala 262:58]
  wire [7:0] combiner_level1_io_s_axis_tkeep_lo = {_combiner_level1_io_s_axis_tkeep_T_23,
    _combiner_level1_io_s_axis_tkeep_T_22,_combiner_level1_io_s_axis_tkeep_T_21,_combiner_level1_io_s_axis_tkeep_T_20,
    _combiner_level1_io_s_axis_tkeep_T_19,_combiner_level1_io_s_axis_tkeep_T_18,_combiner_level1_io_s_axis_tkeep_T_17,
    _combiner_level1_io_s_axis_tkeep_T_16}; // @[bfs_remote.scala 262:87]
  wire [79:0] _combiner_level1_io_s_axis_tkeep_T_32 = {combiner_level1_io_s_axis_tkeep_hi,
    _combiner_level1_io_s_axis_tkeep_T_31,_combiner_level1_io_s_axis_tkeep_T_30,_combiner_level1_io_s_axis_tkeep_T_29,
    _combiner_level1_io_s_axis_tkeep_T_28,_combiner_level1_io_s_axis_tkeep_T_27,_combiner_level1_io_s_axis_tkeep_T_26,
    _combiner_level1_io_s_axis_tkeep_T_25,_combiner_level1_io_s_axis_tkeep_T_24,combiner_level1_io_s_axis_tkeep_lo}; // @[Cat.scala 30:58]
  wire  _combiner_level1_io_s_axis_tvalid_T_1 = xbar_level0_m_axis_tvalid[0] | io_remote_in_valid; // @[bfs_remote.scala 264:91]
  wire  xbar_level0_io_m_axis_tready_lo = combiner_level1_s_axis_tready[1]; // @[bfs_remote.scala 266:92]
  wire [7:0] xbar_level1_io_m_axis_tready_lo = {io_pe_out_7_ready,io_pe_out_6_ready,io_pe_out_5_ready,io_pe_out_4_ready,
    io_pe_out_3_ready,io_pe_out_2_ready,io_pe_out_1_ready,io_pe_out_0_ready}; // @[bfs_remote.scala 280:12]
  wire [7:0] xbar_level1_io_m_axis_tready_hi = {io_pe_out_15_ready,io_pe_out_14_ready,io_pe_out_13_ready,
    io_pe_out_12_ready,io_pe_out_11_ready,io_pe_out_10_ready,io_pe_out_9_ready,io_pe_out_8_ready}; // @[bfs_remote.scala 280:12]
  axis_combiner_level0 combiner_level0 ( // @[bfs_remote.scala 238:31]
    .aclk(combiner_level0_aclk),
    .aresetn(combiner_level0_aresetn),
    .s_axis_tdata(combiner_level0_s_axis_tdata),
    .s_axis_tkeep(combiner_level0_s_axis_tkeep),
    .s_axis_tlast(combiner_level0_s_axis_tlast),
    .s_axis_tvalid(combiner_level0_s_axis_tvalid),
    .s_axis_tready(combiner_level0_s_axis_tready),
    .s_axis_tid(combiner_level0_s_axis_tid),
    .m_axis_tdata(combiner_level0_m_axis_tdata),
    .m_axis_tkeep(combiner_level0_m_axis_tkeep),
    .m_axis_tlast(combiner_level0_m_axis_tlast),
    .m_axis_tvalid(combiner_level0_m_axis_tvalid),
    .m_axis_tready(combiner_level0_m_axis_tready),
    .m_axis_tid(combiner_level0_m_axis_tid)
  );
  axis_broadcaster_level0 xbar_level0 ( // @[bfs_remote.scala 250:27]
    .aclk(xbar_level0_aclk),
    .aresetn(xbar_level0_aresetn),
    .s_axis_tdata(xbar_level0_s_axis_tdata),
    .s_axis_tkeep(xbar_level0_s_axis_tkeep),
    .s_axis_tlast(xbar_level0_s_axis_tlast),
    .s_axis_tvalid(xbar_level0_s_axis_tvalid),
    .s_axis_tready(xbar_level0_s_axis_tready),
    .s_axis_tid(xbar_level0_s_axis_tid),
    .m_axis_tdata(xbar_level0_m_axis_tdata),
    .m_axis_tkeep(xbar_level0_m_axis_tkeep),
    .m_axis_tlast(xbar_level0_m_axis_tlast),
    .m_axis_tvalid(xbar_level0_m_axis_tvalid),
    .m_axis_tready(xbar_level0_m_axis_tready),
    .m_axis_tid(xbar_level0_m_axis_tid)
  );
  axis_combiner_level1 combiner_level1 ( // @[bfs_remote.scala 257:31]
    .aclk(combiner_level1_aclk),
    .aresetn(combiner_level1_aresetn),
    .s_axis_tdata(combiner_level1_s_axis_tdata),
    .s_axis_tkeep(combiner_level1_s_axis_tkeep),
    .s_axis_tlast(combiner_level1_s_axis_tlast),
    .s_axis_tvalid(combiner_level1_s_axis_tvalid),
    .s_axis_tready(combiner_level1_s_axis_tready),
    .s_axis_tid(combiner_level1_s_axis_tid),
    .m_axis_tdata(combiner_level1_m_axis_tdata),
    .m_axis_tkeep(combiner_level1_m_axis_tkeep),
    .m_axis_tlast(combiner_level1_m_axis_tlast),
    .m_axis_tvalid(combiner_level1_m_axis_tvalid),
    .m_axis_tready(combiner_level1_m_axis_tready),
    .m_axis_tid(combiner_level1_m_axis_tid)
  );
  axis_broadcaster_level1 xbar_level1 ( // @[bfs_remote.scala 268:27]
    .aclk(xbar_level1_aclk),
    .aresetn(xbar_level1_aresetn),
    .s_axis_tdata(xbar_level1_s_axis_tdata),
    .s_axis_tkeep(xbar_level1_s_axis_tkeep),
    .s_axis_tlast(xbar_level1_s_axis_tlast),
    .s_axis_tvalid(xbar_level1_s_axis_tvalid),
    .s_axis_tready(xbar_level1_s_axis_tready),
    .s_axis_tid(xbar_level1_s_axis_tid),
    .m_axis_tdata(xbar_level1_m_axis_tdata),
    .m_axis_tkeep(xbar_level1_m_axis_tkeep),
    .m_axis_tlast(xbar_level1_m_axis_tlast),
    .m_axis_tvalid(xbar_level1_m_axis_tvalid),
    .m_axis_tready(xbar_level1_m_axis_tready),
    .m_axis_tid(xbar_level1_m_axis_tid)
  );
  assign io_ddr_in_0_ready = combiner_level0_s_axis_tready[0]; // @[bfs_remote.scala 247:65]
  assign io_ddr_in_1_ready = combiner_level0_s_axis_tready[1]; // @[bfs_remote.scala 247:65]
  assign io_ddr_in_2_ready = combiner_level0_s_axis_tready[2]; // @[bfs_remote.scala 247:65]
  assign io_ddr_in_3_ready = combiner_level0_s_axis_tready[3]; // @[bfs_remote.scala 247:65]
  assign io_pe_out_0_valid = xbar_level1_m_axis_tvalid[0]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_0_bits_tdata = xbar_level1_m_axis_tdata[1023:0]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_0_bits_tkeep = xbar_level1_m_axis_tkeep[31:0]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_1_valid = xbar_level1_m_axis_tvalid[1]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_1_bits_tdata = xbar_level1_m_axis_tdata[2047:1024]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_1_bits_tkeep = xbar_level1_m_axis_tkeep[159:128]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_2_valid = xbar_level1_m_axis_tvalid[2]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_2_bits_tdata = xbar_level1_m_axis_tdata[3071:2048]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_2_bits_tkeep = xbar_level1_m_axis_tkeep[287:256]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_3_valid = xbar_level1_m_axis_tvalid[3]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_3_bits_tdata = xbar_level1_m_axis_tdata[4095:3072]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_3_bits_tkeep = xbar_level1_m_axis_tkeep[415:384]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_4_valid = xbar_level1_m_axis_tvalid[4]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_4_bits_tdata = xbar_level1_m_axis_tdata[5119:4096]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_4_bits_tkeep = xbar_level1_m_axis_tkeep[543:512]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_5_valid = xbar_level1_m_axis_tvalid[5]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_5_bits_tdata = xbar_level1_m_axis_tdata[6143:5120]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_5_bits_tkeep = xbar_level1_m_axis_tkeep[671:640]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_6_valid = xbar_level1_m_axis_tvalid[6]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_6_bits_tdata = xbar_level1_m_axis_tdata[7167:6144]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_6_bits_tkeep = xbar_level1_m_axis_tkeep[799:768]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_7_valid = xbar_level1_m_axis_tvalid[7]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_7_bits_tdata = xbar_level1_m_axis_tdata[8191:7168]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_7_bits_tkeep = xbar_level1_m_axis_tkeep[927:896]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_8_valid = xbar_level1_m_axis_tvalid[8]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_8_bits_tdata = xbar_level1_m_axis_tdata[9215:8192]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_8_bits_tkeep = xbar_level1_m_axis_tkeep[1055:1024]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_9_valid = xbar_level1_m_axis_tvalid[9]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_9_bits_tdata = xbar_level1_m_axis_tdata[10239:9216]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_9_bits_tkeep = xbar_level1_m_axis_tkeep[1183:1152]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_10_valid = xbar_level1_m_axis_tvalid[10]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_10_bits_tdata = xbar_level1_m_axis_tdata[11263:10240]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_10_bits_tkeep = xbar_level1_m_axis_tkeep[1311:1280]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_11_valid = xbar_level1_m_axis_tvalid[11]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_11_bits_tdata = xbar_level1_m_axis_tdata[12287:11264]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_11_bits_tkeep = xbar_level1_m_axis_tkeep[1439:1408]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_12_valid = xbar_level1_m_axis_tvalid[12]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_12_bits_tdata = xbar_level1_m_axis_tdata[13311:12288]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_12_bits_tkeep = xbar_level1_m_axis_tkeep[1567:1536]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_13_valid = xbar_level1_m_axis_tvalid[13]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_13_bits_tdata = xbar_level1_m_axis_tdata[14335:13312]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_13_bits_tkeep = xbar_level1_m_axis_tkeep[1695:1664]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_14_valid = xbar_level1_m_axis_tvalid[14]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_14_bits_tdata = xbar_level1_m_axis_tdata[15359:14336]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_14_bits_tkeep = xbar_level1_m_axis_tkeep[1823:1792]; // @[nf_arm_doce_top.scala 124:13]
  assign io_pe_out_15_valid = xbar_level1_m_axis_tvalid[15]; // @[bfs_remote.scala 275:47]
  assign io_pe_out_15_bits_tdata = xbar_level1_m_axis_tdata[16383:15360]; // @[nf_arm_doce_top.scala 122:21]
  assign io_pe_out_15_bits_tkeep = xbar_level1_m_axis_tkeep[1951:1920]; // @[nf_arm_doce_top.scala 124:13]
  assign io_remote_out_valid = xbar_level0_m_axis_tvalid[1]; // @[bfs_remote.scala 255:54]
  assign io_remote_out_bits_tdata = xbar_level0_m_axis_tdata[1023:512]; // @[nf_arm_doce_top.scala 122:21]
  assign io_remote_out_bits_tkeep = xbar_level0_m_axis_tkeep[79:64]; // @[nf_arm_doce_top.scala 124:13]
  assign io_remote_in_ready = combiner_level1_s_axis_tready[0]; // @[bfs_remote.scala 265:57]
  assign combiner_level0_aclk = clock; // @[bfs_remote.scala 239:42]
  assign combiner_level0_aresetn = ~reset; // @[bfs_remote.scala 240:33]
  assign combiner_level0_s_axis_tdata = {combiner_level0_io_s_axis_tdata_hi,combiner_level0_io_s_axis_tdata_lo}; // @[bfs_remote.scala 241:103]
  assign combiner_level0_s_axis_tkeep = {{48'd0}, _combiner_level0_io_s_axis_tkeep_T_32}; // @[bfs_remote.scala 243:33]
  assign combiner_level0_s_axis_tlast = 4'hf; // @[bfs_remote.scala 244:103]
  assign combiner_level0_s_axis_tvalid = {combiner_level0_io_s_axis_tvalid_lo,combiner_level0_io_s_axis_tvalid_lo}; // @[bfs_remote.scala 245:116]
  assign combiner_level0_s_axis_tid = 4'h0;
  assign combiner_level0_m_axis_tready = xbar_level0_s_axis_tready; // @[bfs_remote.scala 253:25]
  assign xbar_level0_aclk = clock; // @[bfs_remote.scala 251:38]
  assign xbar_level0_aresetn = ~reset; // @[bfs_remote.scala 252:29]
  assign xbar_level0_s_axis_tdata = combiner_level0_m_axis_tdata; // @[bfs_remote.scala 253:25]
  assign xbar_level0_s_axis_tkeep = combiner_level0_m_axis_tkeep; // @[bfs_remote.scala 253:25]
  assign xbar_level0_s_axis_tlast = combiner_level0_m_axis_tlast; // @[bfs_remote.scala 253:25]
  assign xbar_level0_s_axis_tvalid = combiner_level0_m_axis_tvalid; // @[bfs_remote.scala 253:25]
  assign xbar_level0_s_axis_tid = combiner_level0_m_axis_tid; // @[bfs_remote.scala 253:25]
  assign xbar_level0_m_axis_tready = {io_remote_out_ready,xbar_level0_io_m_axis_tready_lo}; // @[Cat.scala 30:58]
  assign combiner_level1_aclk = clock; // @[bfs_remote.scala 258:42]
  assign combiner_level1_aresetn = ~reset; // @[bfs_remote.scala 259:33]
  assign combiner_level1_s_axis_tdata = {combiner_level1_io_s_axis_tdata_hi,io_remote_in_bits_tdata}; // @[Cat.scala 30:58]
  assign combiner_level1_s_axis_tkeep = {{48'd0}, _combiner_level1_io_s_axis_tkeep_T_32}; // @[Cat.scala 30:58]
  assign combiner_level1_s_axis_tlast = 2'h3; // @[bfs_remote.scala 263:35]
  assign combiner_level1_s_axis_tvalid = {_combiner_level1_io_s_axis_tvalid_T_1,_combiner_level1_io_s_axis_tvalid_T_1}; // @[bfs_remote.scala 264:120]
  assign combiner_level1_s_axis_tid = 2'h0;
  assign combiner_level1_m_axis_tready = xbar_level1_s_axis_tready; // @[bfs_remote.scala 271:25]
  assign xbar_level1_aclk = clock; // @[bfs_remote.scala 269:38]
  assign xbar_level1_aresetn = ~reset; // @[bfs_remote.scala 270:29]
  assign xbar_level1_s_axis_tdata = combiner_level1_m_axis_tdata; // @[bfs_remote.scala 271:25]
  assign xbar_level1_s_axis_tkeep = combiner_level1_m_axis_tkeep; // @[bfs_remote.scala 271:25]
  assign xbar_level1_s_axis_tlast = combiner_level1_m_axis_tlast; // @[bfs_remote.scala 271:25]
  assign xbar_level1_s_axis_tvalid = combiner_level1_m_axis_tvalid; // @[bfs_remote.scala 271:25]
  assign xbar_level1_s_axis_tid = combiner_level1_m_axis_tid; // @[bfs_remote.scala 271:25]
  assign xbar_level1_m_axis_tready = {xbar_level1_io_m_axis_tready_hi,xbar_level1_io_m_axis_tready_lo}; // @[bfs_remote.scala 280:12]
endmodule
module Remote_Apply(
  input          clock,
  input          reset,
  output         io_xbar_in_ready,
  input          io_xbar_in_valid,
  input  [511:0] io_xbar_in_bits_tdata,
  input  [15:0]  io_xbar_in_bits_tkeep,
  input          io_remote_out_aw_ready,
  output         io_remote_out_aw_valid,
  output [63:0]  io_remote_out_aw_bits_awaddr,
  output [5:0]   io_remote_out_aw_bits_awid,
  input          io_remote_out_w_ready,
  output         io_remote_out_w_valid,
  output [511:0] io_remote_out_w_bits_wdata,
  output [63:0]  io_remote_out_w_bits_wstrb,
  input  [3:0]   io_recv_sync,
  input          io_recv_sync_phase2,
  input          io_signal,
  output         io_signal_ack,
  input          io_local_fpga_id,
  input  [63:0]  io_level_base_addr,
  input  [31:0]  io_local_unvisited_size,
  output         io_end
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_in_fifo_s_axis_aclk; // @[bfs_remote.scala 54:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[bfs_remote.scala 54:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[bfs_remote.scala 54:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[bfs_remote.scala 54:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[bfs_remote.scala 54:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[bfs_remote.scala 54:30]
  wire  vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 54:30]
  wire  vertex_in_fifo_s_axis_tid; // @[bfs_remote.scala 54:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 54:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 54:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[bfs_remote.scala 54:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 54:30]
  wire  vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 54:30]
  wire  vertex_in_fifo_m_axis_tid; // @[bfs_remote.scala 54:30]
  wire  _filtered_keep_0_T_5 = io_xbar_in_bits_tdata[4] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_0_T_6 = io_xbar_in_bits_tdata[31] ? 1'h0 : _filtered_keep_0_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_0 = io_xbar_in_bits_tkeep[0] & _filtered_keep_0_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_1_T_5 = io_xbar_in_bits_tdata[36] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_1_T_6 = io_xbar_in_bits_tdata[63] ? 1'h0 : _filtered_keep_1_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_1 = io_xbar_in_bits_tkeep[1] & _filtered_keep_1_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_2_T_5 = io_xbar_in_bits_tdata[68] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_2_T_6 = io_xbar_in_bits_tdata[95] ? 1'h0 : _filtered_keep_2_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_2 = io_xbar_in_bits_tkeep[2] & _filtered_keep_2_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_3_T_5 = io_xbar_in_bits_tdata[100] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_3_T_6 = io_xbar_in_bits_tdata[127] ? 1'h0 : _filtered_keep_3_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_3 = io_xbar_in_bits_tkeep[3] & _filtered_keep_3_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_4_T_5 = io_xbar_in_bits_tdata[132] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_4_T_6 = io_xbar_in_bits_tdata[159] ? 1'h0 : _filtered_keep_4_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_4 = io_xbar_in_bits_tkeep[4] & _filtered_keep_4_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_5_T_5 = io_xbar_in_bits_tdata[164] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_5_T_6 = io_xbar_in_bits_tdata[191] ? 1'h0 : _filtered_keep_5_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_5 = io_xbar_in_bits_tkeep[5] & _filtered_keep_5_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_6_T_5 = io_xbar_in_bits_tdata[196] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_6_T_6 = io_xbar_in_bits_tdata[223] ? 1'h0 : _filtered_keep_6_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_6 = io_xbar_in_bits_tkeep[6] & _filtered_keep_6_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_7_T_5 = io_xbar_in_bits_tdata[228] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_7_T_6 = io_xbar_in_bits_tdata[255] ? 1'h0 : _filtered_keep_7_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_7 = io_xbar_in_bits_tkeep[7] & _filtered_keep_7_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_8_T_5 = io_xbar_in_bits_tdata[260] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_8_T_6 = io_xbar_in_bits_tdata[287] ? 1'h0 : _filtered_keep_8_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_8 = io_xbar_in_bits_tkeep[8] & _filtered_keep_8_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_9_T_5 = io_xbar_in_bits_tdata[292] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_9_T_6 = io_xbar_in_bits_tdata[319] ? 1'h0 : _filtered_keep_9_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_9 = io_xbar_in_bits_tkeep[9] & _filtered_keep_9_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_10_T_5 = io_xbar_in_bits_tdata[324] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_10_T_6 = io_xbar_in_bits_tdata[351] ? 1'h0 : _filtered_keep_10_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_10 = io_xbar_in_bits_tkeep[10] & _filtered_keep_10_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_11_T_5 = io_xbar_in_bits_tdata[356] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_11_T_6 = io_xbar_in_bits_tdata[383] ? 1'h0 : _filtered_keep_11_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_11 = io_xbar_in_bits_tkeep[11] & _filtered_keep_11_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_12_T_5 = io_xbar_in_bits_tdata[388] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_12_T_6 = io_xbar_in_bits_tdata[415] ? 1'h0 : _filtered_keep_12_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_12 = io_xbar_in_bits_tkeep[12] & _filtered_keep_12_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_13_T_5 = io_xbar_in_bits_tdata[420] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_13_T_6 = io_xbar_in_bits_tdata[447] ? 1'h0 : _filtered_keep_13_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_13 = io_xbar_in_bits_tkeep[13] & _filtered_keep_13_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_14_T_5 = io_xbar_in_bits_tdata[452] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_14_T_6 = io_xbar_in_bits_tdata[479] ? 1'h0 : _filtered_keep_14_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_14 = io_xbar_in_bits_tkeep[14] & _filtered_keep_14_T_6; // @[bfs_remote.scala 48:15]
  wire  _filtered_keep_15_T_5 = io_xbar_in_bits_tdata[484] != io_local_fpga_id; // @[bfs_remote.scala 35:88]
  wire  _filtered_keep_15_T_6 = io_xbar_in_bits_tdata[511] ? 1'h0 : _filtered_keep_15_T_5; // @[bfs_remote.scala 49:12]
  wire  filtered_keep_15 = io_xbar_in_bits_tkeep[15] & _filtered_keep_15_T_6; // @[bfs_remote.scala 48:15]
  wire [63:0] _GEN_29 = {{32'd0}, io_local_unvisited_size}; // @[bfs_remote.scala 65:57]
  wire [63:0] sync_data = 64'h80000000 + _GEN_29; // @[bfs_remote.scala 65:57]
  (*dont_touch = "true" *)reg [2:0] sync_status; // @[bfs_remote.scala 66:28]
  wire  _T_3 = sync_status == 3'h4; // @[bfs_remote.scala 69:26]
  wire  _T_4 = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 69:92]
  wire  _T_8 = sync_status == 3'h6; // @[bfs_remote.scala 73:26]
  wire [2:0] _GEN_0 = sync_status == 3'h7 & io_signal ? 3'h0 : sync_status; // @[bfs_remote.scala 75:58 bfs_remote.scala 76:17 bfs_remote.scala 66:28]
  wire [2:0] _GEN_1 = sync_status == 3'h6 & _T_4 ? 3'h7 : _GEN_0; // @[bfs_remote.scala 73:95 bfs_remote.scala 74:17]
  wire  need_to_send_sync = _T_3 | _T_8; // @[bfs_remote.scala 80:66]
  wire [7:0] vertex_in_fifo_io_s_axis_tkeep_lo = {filtered_keep_7,filtered_keep_6,filtered_keep_5,filtered_keep_4,
    filtered_keep_3,filtered_keep_2,filtered_keep_1,filtered_keep_0}; // @[bfs_remote.scala 85:85]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T = {filtered_keep_15,filtered_keep_14,filtered_keep_13,filtered_keep_12,
    filtered_keep_11,filtered_keep_10,filtered_keep_9,filtered_keep_8,vertex_in_fifo_io_s_axis_tkeep_lo}; // @[bfs_remote.scala 85:85]
  wire [15:0] _vertex_in_fifo_io_s_axis_tkeep_T_1 = need_to_send_sync ? 16'h1 : _vertex_in_fifo_io_s_axis_tkeep_T; // @[bfs_remote.scala 85:40]
  reg [2:0] send_status; // @[bfs_remote.scala 92:28]
  wire [511:0] _dest_next_WIRE_1 = vertex_in_fifo_m_axis_tdata;
  wire  _dest_next_T_37 = ~_dest_next_WIRE_1[4] | _dest_next_WIRE_1[31]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_40 = _dest_next_T_37 & vertex_in_fifo_m_axis_tkeep[0] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_45 = ~_dest_next_WIRE_1[36] | _dest_next_WIRE_1[63]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_48 = _dest_next_T_45 & vertex_in_fifo_m_axis_tkeep[1] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_53 = ~_dest_next_WIRE_1[68] | _dest_next_WIRE_1[95]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_56 = _dest_next_T_53 & vertex_in_fifo_m_axis_tkeep[2] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_61 = ~_dest_next_WIRE_1[100] | _dest_next_WIRE_1[127]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_64 = _dest_next_T_61 & vertex_in_fifo_m_axis_tkeep[3] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_69 = ~_dest_next_WIRE_1[132] | _dest_next_WIRE_1[159]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_72 = _dest_next_T_69 & vertex_in_fifo_m_axis_tkeep[4] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_77 = ~_dest_next_WIRE_1[164] | _dest_next_WIRE_1[191]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_80 = _dest_next_T_77 & vertex_in_fifo_m_axis_tkeep[5] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_85 = ~_dest_next_WIRE_1[196] | _dest_next_WIRE_1[223]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_88 = _dest_next_T_85 & vertex_in_fifo_m_axis_tkeep[6] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_93 = ~_dest_next_WIRE_1[228] | _dest_next_WIRE_1[255]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_96 = _dest_next_T_93 & vertex_in_fifo_m_axis_tkeep[7] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_101 = ~_dest_next_WIRE_1[260] | _dest_next_WIRE_1[287]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_104 = _dest_next_T_101 & vertex_in_fifo_m_axis_tkeep[8] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_109 = ~_dest_next_WIRE_1[292] | _dest_next_WIRE_1[319]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_112 = _dest_next_T_109 & vertex_in_fifo_m_axis_tkeep[9] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_117 = ~_dest_next_WIRE_1[324] | _dest_next_WIRE_1[351]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_120 = _dest_next_T_117 & vertex_in_fifo_m_axis_tkeep[10] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_125 = ~_dest_next_WIRE_1[356] | _dest_next_WIRE_1[383]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_128 = _dest_next_T_125 & vertex_in_fifo_m_axis_tkeep[11] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_133 = ~_dest_next_WIRE_1[388] | _dest_next_WIRE_1[415]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_136 = _dest_next_T_133 & vertex_in_fifo_m_axis_tkeep[12] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_141 = ~_dest_next_WIRE_1[420] | _dest_next_WIRE_1[447]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_144 = _dest_next_T_141 & vertex_in_fifo_m_axis_tkeep[13] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_149 = ~_dest_next_WIRE_1[452] | _dest_next_WIRE_1[479]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_152 = _dest_next_T_149 & vertex_in_fifo_m_axis_tkeep[14] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_157 = ~_dest_next_WIRE_1[484] | _dest_next_WIRE_1[511]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_160 = _dest_next_T_157 & vertex_in_fifo_m_axis_tkeep[15] & io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  dest_next_0 = _dest_next_T_40 | _dest_next_T_48 | _dest_next_T_56 | _dest_next_T_64 | _dest_next_T_72 |
    _dest_next_T_80 | _dest_next_T_88 | _dest_next_T_96 | _dest_next_T_104 | _dest_next_T_112 | _dest_next_T_120 |
    _dest_next_T_128 | _dest_next_T_136 | _dest_next_T_144 | _dest_next_T_152 | _dest_next_T_160; // @[bfs_remote.scala 95:85]
  wire  _dest_next_T_213 = _dest_next_WIRE_1[4] | _dest_next_WIRE_1[31]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_216 = _dest_next_T_213 & vertex_in_fifo_m_axis_tkeep[0] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_221 = _dest_next_WIRE_1[36] | _dest_next_WIRE_1[63]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_224 = _dest_next_T_221 & vertex_in_fifo_m_axis_tkeep[1] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_229 = _dest_next_WIRE_1[68] | _dest_next_WIRE_1[95]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_232 = _dest_next_T_229 & vertex_in_fifo_m_axis_tkeep[2] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_237 = _dest_next_WIRE_1[100] | _dest_next_WIRE_1[127]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_240 = _dest_next_T_237 & vertex_in_fifo_m_axis_tkeep[3] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_245 = _dest_next_WIRE_1[132] | _dest_next_WIRE_1[159]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_248 = _dest_next_T_245 & vertex_in_fifo_m_axis_tkeep[4] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_253 = _dest_next_WIRE_1[164] | _dest_next_WIRE_1[191]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_256 = _dest_next_T_253 & vertex_in_fifo_m_axis_tkeep[5] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_261 = _dest_next_WIRE_1[196] | _dest_next_WIRE_1[223]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_264 = _dest_next_T_261 & vertex_in_fifo_m_axis_tkeep[6] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_269 = _dest_next_WIRE_1[228] | _dest_next_WIRE_1[255]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_272 = _dest_next_T_269 & vertex_in_fifo_m_axis_tkeep[7] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_277 = _dest_next_WIRE_1[260] | _dest_next_WIRE_1[287]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_280 = _dest_next_T_277 & vertex_in_fifo_m_axis_tkeep[8] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_285 = _dest_next_WIRE_1[292] | _dest_next_WIRE_1[319]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_288 = _dest_next_T_285 & vertex_in_fifo_m_axis_tkeep[9] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_293 = _dest_next_WIRE_1[324] | _dest_next_WIRE_1[351]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_296 = _dest_next_T_293 & vertex_in_fifo_m_axis_tkeep[10] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_301 = _dest_next_WIRE_1[356] | _dest_next_WIRE_1[383]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_304 = _dest_next_T_301 & vertex_in_fifo_m_axis_tkeep[11] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_309 = _dest_next_WIRE_1[388] | _dest_next_WIRE_1[415]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_312 = _dest_next_T_309 & vertex_in_fifo_m_axis_tkeep[12] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_317 = _dest_next_WIRE_1[420] | _dest_next_WIRE_1[447]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_320 = _dest_next_T_317 & vertex_in_fifo_m_axis_tkeep[13] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_325 = _dest_next_WIRE_1[452] | _dest_next_WIRE_1[479]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_328 = _dest_next_T_325 & vertex_in_fifo_m_axis_tkeep[14] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _dest_next_T_333 = _dest_next_WIRE_1[484] | _dest_next_WIRE_1[511]; // @[bfs_remote.scala 40:116]
  wire  _dest_next_T_336 = _dest_next_T_333 & vertex_in_fifo_m_axis_tkeep[15] & ~io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  dest_next_1 = _dest_next_T_216 | _dest_next_T_224 | _dest_next_T_232 | _dest_next_T_240 | _dest_next_T_248 |
    _dest_next_T_256 | _dest_next_T_264 | _dest_next_T_272 | _dest_next_T_280 | _dest_next_T_288 | _dest_next_T_296 |
    _dest_next_T_304 | _dest_next_T_312 | _dest_next_T_320 | _dest_next_T_328 | _dest_next_T_336; // @[bfs_remote.scala 95:85]
  reg  dest_0; // @[bfs_remote.scala 97:21]
  reg [31:0] count; // @[bfs_remote.scala 99:22]
  wire  last_send = send_status != 3'h0 & count == 32'h1; // @[bfs_remote.scala 100:44]
  wire  addr_issue = io_remote_out_aw_valid & io_remote_out_aw_ready; // @[bfs_remote.scala 101:43]
  wire  data_issue = io_remote_out_w_valid & io_remote_out_w_ready; // @[bfs_remote.scala 102:42]
  wire  dest_grant = dest_0 ? 1'h0 : 1'h1; // @[bfs_remote.scala 105:18 bfs_remote.scala 106:18 bfs_remote.scala 103:14]
  wire [31:0] _count_WIRE = {{31'd0}, dest_next_0}; // @[bfs_remote.scala 114:45 bfs_remote.scala 114:45]
  wire [31:0] _count_WIRE_1 = {{31'd0}, dest_next_1}; // @[bfs_remote.scala 114:45 bfs_remote.scala 114:45]
  wire [31:0] _count_T_1 = _count_WIRE + _count_WIRE_1; // @[bfs_remote.scala 114:67]
  wire  _GEN_10 = dest_next_0 | dest_next_1 ? 1'h0 : 1'h1; // @[bfs_remote.scala 111:33 bfs_remote.scala 109:35 bfs_remote.scala 116:39]
  wire  _T_17 = send_status == 3'h1; // @[bfs_remote.scala 118:27]
  wire  _T_18 = send_status == 3'h1 & addr_issue; // @[bfs_remote.scala 118:42]
  wire  _T_19 = send_status == 3'h1 & addr_issue & data_issue; // @[bfs_remote.scala 118:56]
  wire  _T_20 = send_status == 3'h2; // @[bfs_remote.scala 119:19]
  wire  _T_22 = _T_19 | send_status == 3'h2 & addr_issue; // @[bfs_remote.scala 119:3]
  wire  _T_23 = send_status == 3'h3; // @[bfs_remote.scala 120:19]
  wire  _dest_0_T_1 = ~dest_grant ? 1'h0 : dest_0; // @[bfs_remote.scala 128:19]
  wire [31:0] _count_T_3 = count - 32'h1; // @[bfs_remote.scala 131:22]
  wire [2:0] _GEN_16 = _T_18 & ~data_issue ? 3'h3 : send_status; // @[bfs_remote.scala 135:70 bfs_remote.scala 136:17 bfs_remote.scala 92:28]
  wire  _GEN_20 = (_T_22 | send_status == 3'h3 & data_issue) & last_send; // @[bfs_remote.scala 120:48 bfs_remote.scala 109:35]
  wire  _io_remote_out_w_bits_wstrb_T_37 = _dest_next_WIRE_1[4] == dest_grant | _dest_next_WIRE_1[31]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_40 = _io_remote_out_w_bits_wstrb_T_37 & vertex_in_fifo_m_axis_tkeep[0] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_45 = _dest_next_WIRE_1[36] == dest_grant | _dest_next_WIRE_1[63]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_48 = _io_remote_out_w_bits_wstrb_T_45 & vertex_in_fifo_m_axis_tkeep[1] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_53 = _dest_next_WIRE_1[68] == dest_grant | _dest_next_WIRE_1[95]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_56 = _io_remote_out_w_bits_wstrb_T_53 & vertex_in_fifo_m_axis_tkeep[2] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_61 = _dest_next_WIRE_1[100] == dest_grant | _dest_next_WIRE_1[127]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_64 = _io_remote_out_w_bits_wstrb_T_61 & vertex_in_fifo_m_axis_tkeep[3] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_69 = _dest_next_WIRE_1[132] == dest_grant | _dest_next_WIRE_1[159]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_72 = _io_remote_out_w_bits_wstrb_T_69 & vertex_in_fifo_m_axis_tkeep[4] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_77 = _dest_next_WIRE_1[164] == dest_grant | _dest_next_WIRE_1[191]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_80 = _io_remote_out_w_bits_wstrb_T_77 & vertex_in_fifo_m_axis_tkeep[5] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_85 = _dest_next_WIRE_1[196] == dest_grant | _dest_next_WIRE_1[223]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_88 = _io_remote_out_w_bits_wstrb_T_85 & vertex_in_fifo_m_axis_tkeep[6] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_93 = _dest_next_WIRE_1[228] == dest_grant | _dest_next_WIRE_1[255]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_96 = _io_remote_out_w_bits_wstrb_T_93 & vertex_in_fifo_m_axis_tkeep[7] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_101 = _dest_next_WIRE_1[260] == dest_grant | _dest_next_WIRE_1[287]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_104 = _io_remote_out_w_bits_wstrb_T_101 & vertex_in_fifo_m_axis_tkeep[8] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_109 = _dest_next_WIRE_1[292] == dest_grant | _dest_next_WIRE_1[319]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_112 = _io_remote_out_w_bits_wstrb_T_109 & vertex_in_fifo_m_axis_tkeep[9] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_117 = _dest_next_WIRE_1[324] == dest_grant | _dest_next_WIRE_1[351]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_120 = _io_remote_out_w_bits_wstrb_T_117 & vertex_in_fifo_m_axis_tkeep[10] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_125 = _dest_next_WIRE_1[356] == dest_grant | _dest_next_WIRE_1[383]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_128 = _io_remote_out_w_bits_wstrb_T_125 & vertex_in_fifo_m_axis_tkeep[11] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_133 = _dest_next_WIRE_1[388] == dest_grant | _dest_next_WIRE_1[415]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_136 = _io_remote_out_w_bits_wstrb_T_133 & vertex_in_fifo_m_axis_tkeep[12] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_141 = _dest_next_WIRE_1[420] == dest_grant | _dest_next_WIRE_1[447]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_144 = _io_remote_out_w_bits_wstrb_T_141 & vertex_in_fifo_m_axis_tkeep[13] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_149 = _dest_next_WIRE_1[452] == dest_grant | _dest_next_WIRE_1[479]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_152 = _io_remote_out_w_bits_wstrb_T_149 & vertex_in_fifo_m_axis_tkeep[14] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire  _io_remote_out_w_bits_wstrb_T_157 = _dest_next_WIRE_1[484] == dest_grant | _dest_next_WIRE_1[511]; // @[bfs_remote.scala 40:116]
  wire  _io_remote_out_w_bits_wstrb_T_160 = _io_remote_out_w_bits_wstrb_T_157 & vertex_in_fifo_m_axis_tkeep[15] &
    dest_grant != io_local_fpga_id; // @[bfs_remote.scala 41:50]
  wire [7:0] io_remote_out_w_bits_wstrb_lo = {_io_remote_out_w_bits_wstrb_T_96,_io_remote_out_w_bits_wstrb_T_88,
    _io_remote_out_w_bits_wstrb_T_80,_io_remote_out_w_bits_wstrb_T_72,_io_remote_out_w_bits_wstrb_T_64,
    _io_remote_out_w_bits_wstrb_T_56,_io_remote_out_w_bits_wstrb_T_48,_io_remote_out_w_bits_wstrb_T_40}; // @[bfs_remote.scala 153:94]
  wire [15:0] _io_remote_out_w_bits_wstrb_T_161 = {_io_remote_out_w_bits_wstrb_T_160,_io_remote_out_w_bits_wstrb_T_152,
    _io_remote_out_w_bits_wstrb_T_144,_io_remote_out_w_bits_wstrb_T_136,_io_remote_out_w_bits_wstrb_T_128,
    _io_remote_out_w_bits_wstrb_T_120,_io_remote_out_w_bits_wstrb_T_112,_io_remote_out_w_bits_wstrb_T_104,
    io_remote_out_w_bits_wstrb_lo}; // @[bfs_remote.scala 153:94]
  (*dont_touch = "true" *)reg [31:0] packet_sent; // @[bfs_remote.scala 155:28]
  wire [31:0] _packet_sent_T_1 = packet_sent + 32'h1; // @[bfs_remote.scala 158:32]
  remote_vid_fifo vertex_in_fifo ( // @[bfs_remote.scala 54:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  assign io_xbar_in_ready = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 88:20]
  assign io_remote_out_aw_valid = _T_17 | _T_20; // @[bfs_remote.scala 140:56]
  assign io_remote_out_aw_bits_awaddr = io_level_base_addr; // @[bfs_remote.scala 146:32]
  assign io_remote_out_aw_bits_awid = {{5'd0}, dest_grant}; // @[bfs_remote.scala 105:18 bfs_remote.scala 106:18 bfs_remote.scala 103:14]
  assign io_remote_out_w_valid = _T_17 | _T_23; // @[bfs_remote.scala 149:55]
  assign io_remote_out_w_bits_wdata = vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 151:30]
  assign io_remote_out_w_bits_wstrb = {{48'd0}, _io_remote_out_w_bits_wstrb_T_161}; // @[bfs_remote.scala 153:94]
  assign io_signal_ack = sync_status == 3'h7; // @[bfs_remote.scala 78:32]
  assign io_end = _T_8 & _T_4; // @[bfs_remote.scala 89:50]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[bfs_remote.scala 81:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[bfs_remote.scala 82:39]
  assign vertex_in_fifo_s_axis_tdata = need_to_send_sync ? {{448'd0}, sync_data} : io_xbar_in_bits_tdata; // @[bfs_remote.scala 87:40]
  assign vertex_in_fifo_s_axis_tkeep = {{48'd0}, _vertex_in_fifo_io_s_axis_tkeep_T_1}; // @[bfs_remote.scala 85:40]
  assign vertex_in_fifo_s_axis_tlast = 1'h1; // @[bfs_remote.scala 86:34]
  assign vertex_in_fifo_s_axis_tvalid = io_xbar_in_valid | need_to_send_sync; // @[bfs_remote.scala 83:57]
  assign vertex_in_fifo_s_axis_tid = 1'h0; // @[bfs_remote.scala 84:32]
  assign vertex_in_fifo_m_axis_tready = send_status == 3'h0 & vertex_in_fifo_m_axis_tvalid ? _GEN_10 : _GEN_20; // @[bfs_remote.scala 110:77]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 66:28]
      sync_status <= 3'h0; // @[bfs_remote.scala 66:28]
    end else if (sync_status == 3'h0 & &io_recv_sync) begin // @[bfs_remote.scala 67:57]
      sync_status <= 3'h4; // @[bfs_remote.scala 68:17]
    end else if (sync_status == 3'h4 & vertex_in_fifo_s_axis_tready) begin // @[bfs_remote.scala 69:95]
      sync_status <= 3'h5; // @[bfs_remote.scala 70:17]
    end else if (sync_status == 3'h5 & io_recv_sync_phase2) begin // @[bfs_remote.scala 71:73]
      sync_status <= 3'h6; // @[bfs_remote.scala 72:17]
    end else begin
      sync_status <= _GEN_1;
    end
    if (reset) begin // @[bfs_remote.scala 92:28]
      send_status <= 3'h0; // @[bfs_remote.scala 92:28]
    end else if (send_status == 3'h0 & vertex_in_fifo_m_axis_tvalid) begin // @[bfs_remote.scala 110:77]
      if (dest_next_0 | dest_next_1) begin // @[bfs_remote.scala 111:33]
        send_status <= 3'h1; // @[bfs_remote.scala 113:19]
      end
    end else if (_T_22 | send_status == 3'h3 & data_issue) begin // @[bfs_remote.scala 120:48]
      if (last_send) begin // @[bfs_remote.scala 121:21]
        send_status <= 3'h0; // @[bfs_remote.scala 123:19]
      end
    end else if (_T_17 & ~addr_issue & data_issue) begin // @[bfs_remote.scala 133:70]
      send_status <= 3'h2; // @[bfs_remote.scala 134:17]
    end else begin
      send_status <= _GEN_16;
    end
    if (reset) begin // @[bfs_remote.scala 97:21]
      dest_0 <= 1'h0; // @[bfs_remote.scala 97:21]
    end else if (send_status == 3'h0 & vertex_in_fifo_m_axis_tvalid) begin // @[bfs_remote.scala 110:77]
      if (dest_next_0 | dest_next_1) begin // @[bfs_remote.scala 111:33]
        dest_0 <= dest_next_0; // @[bfs_remote.scala 112:12]
      end
    end else if (_T_22 | send_status == 3'h3 & data_issue) begin // @[bfs_remote.scala 120:48]
      if (!(last_send)) begin // @[bfs_remote.scala 121:21]
        dest_0 <= _dest_0_T_1; // @[bfs_remote.scala 128:13]
      end
    end
    if (reset) begin // @[bfs_remote.scala 99:22]
      count <= 32'h0; // @[bfs_remote.scala 99:22]
    end else if (send_status == 3'h0 & vertex_in_fifo_m_axis_tvalid) begin // @[bfs_remote.scala 110:77]
      if (dest_next_0 | dest_next_1) begin // @[bfs_remote.scala 111:33]
        count <= _count_T_1; // @[bfs_remote.scala 114:13]
      end
    end else if (_T_22 | send_status == 3'h3 & data_issue) begin // @[bfs_remote.scala 120:48]
      if (last_send) begin // @[bfs_remote.scala 121:21]
        count <= 32'h0; // @[bfs_remote.scala 122:13]
      end else begin
        count <= _count_T_3; // @[bfs_remote.scala 131:13]
      end
    end
    if (reset) begin // @[bfs_remote.scala 155:28]
      packet_sent <= 32'h0; // @[bfs_remote.scala 155:28]
    end else if (addr_issue) begin // @[bfs_remote.scala 157:57]
      packet_sent <= _packet_sent_T_1; // @[bfs_remote.scala 158:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_status = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  send_status = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dest_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  packet_sent = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Remote_Scatter(
  input          clock,
  input          reset,
  output         io_remote_in_w_ready,
  input          io_remote_in_w_valid,
  input  [511:0] io_remote_in_w_bits_wdata,
  input  [63:0]  io_remote_in_w_bits_wstrb,
  input          io_xbar_out_ready,
  output         io_xbar_out_valid,
  output [511:0] io_xbar_out_bits_tdata,
  output [15:0]  io_xbar_out_bits_tkeep,
  input          io_signal,
  input          io_start,
  output         io_issue_sync,
  output         io_issue_sync_phase2,
  output [31:0]  io_remote_unvisited_size
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  vertex_in_fifo_s_axis_aclk; // @[bfs_remote.scala 182:30]
  wire  vertex_in_fifo_s_axis_aresetn; // @[bfs_remote.scala 182:30]
  wire [511:0] vertex_in_fifo_s_axis_tdata; // @[bfs_remote.scala 182:30]
  wire [63:0] vertex_in_fifo_s_axis_tkeep; // @[bfs_remote.scala 182:30]
  wire  vertex_in_fifo_s_axis_tlast; // @[bfs_remote.scala 182:30]
  wire  vertex_in_fifo_s_axis_tvalid; // @[bfs_remote.scala 182:30]
  wire  vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 182:30]
  wire  vertex_in_fifo_s_axis_tid; // @[bfs_remote.scala 182:30]
  wire [511:0] vertex_in_fifo_m_axis_tdata; // @[bfs_remote.scala 182:30]
  wire [63:0] vertex_in_fifo_m_axis_tkeep; // @[bfs_remote.scala 182:30]
  wire  vertex_in_fifo_m_axis_tlast; // @[bfs_remote.scala 182:30]
  wire  vertex_in_fifo_m_axis_tvalid; // @[bfs_remote.scala 182:30]
  wire  vertex_in_fifo_m_axis_tready; // @[bfs_remote.scala 182:30]
  wire  vertex_in_fifo_m_axis_tid; // @[bfs_remote.scala 182:30]
  (*dont_touch = "true" *)reg [1:0] sync; // @[bfs_remote.scala 190:21]
  wire  is_sync = vertex_in_fifo_m_axis_tvalid & vertex_in_fifo_m_axis_tdata[31] & vertex_in_fifo_m_axis_tkeep[0]; // @[bfs_remote.scala 191:104]
  wire [1:0] _sync_T_1 = sync + 2'h1; // @[bfs_remote.scala 196:18]
  wire  _T_1 = ~io_start & io_signal; // @[bfs_remote.scala 197:24]
  wire [63:0] _io_xbar_out_bits_tkeep_T = vertex_in_fifo_m_axis_tkeep; // @[nf_arm_doce_top.scala 124:21]
  wire  _vertex_in_fifo_io_m_axis_tready_T = io_issue_sync ? 1'h0 : io_xbar_out_ready; // @[Mux.scala 98:16]
  wire  _io_xbar_out_valid_T = io_issue_sync ? 1'h0 : vertex_in_fifo_m_axis_tvalid; // @[Mux.scala 98:16]
  (*dont_touch = "true" *)reg [31:0] unvisited_size_reg; // @[bfs_remote.scala 210:35]
  wire [31:0] _GEN_5 = {{1'd0}, vertex_in_fifo_m_axis_tdata[30:0]}; // @[bfs_remote.scala 212:46]
  wire [31:0] _unvisited_size_reg_T_2 = unvisited_size_reg + _GEN_5; // @[bfs_remote.scala 212:46]
  (*dont_touch = "true" *)reg [31:0] packet_recv; // @[bfs_remote.scala 221:28]
  wire [31:0] _packet_recv_T_1 = packet_recv + 32'h1; // @[bfs_remote.scala 224:32]
  remote_vid_fifo vertex_in_fifo ( // @[bfs_remote.scala 182:30]
    .s_axis_aclk(vertex_in_fifo_s_axis_aclk),
    .s_axis_aresetn(vertex_in_fifo_s_axis_aresetn),
    .s_axis_tdata(vertex_in_fifo_s_axis_tdata),
    .s_axis_tkeep(vertex_in_fifo_s_axis_tkeep),
    .s_axis_tlast(vertex_in_fifo_s_axis_tlast),
    .s_axis_tvalid(vertex_in_fifo_s_axis_tvalid),
    .s_axis_tready(vertex_in_fifo_s_axis_tready),
    .s_axis_tid(vertex_in_fifo_s_axis_tid),
    .m_axis_tdata(vertex_in_fifo_m_axis_tdata),
    .m_axis_tkeep(vertex_in_fifo_m_axis_tkeep),
    .m_axis_tlast(vertex_in_fifo_m_axis_tlast),
    .m_axis_tvalid(vertex_in_fifo_m_axis_tvalid),
    .m_axis_tready(vertex_in_fifo_m_axis_tready),
    .m_axis_tid(vertex_in_fifo_m_axis_tid)
  );
  assign io_remote_in_w_ready = vertex_in_fifo_s_axis_tready; // @[bfs_remote.scala 188:24]
  assign io_xbar_out_valid = is_sync ? 1'h0 : _io_xbar_out_valid_T; // @[Mux.scala 98:16]
  assign io_xbar_out_bits_tdata = vertex_in_fifo_m_axis_tdata; // @[nf_arm_doce_top.scala 122:21]
  assign io_xbar_out_bits_tkeep = _io_xbar_out_bits_tkeep_T[15:0]; // @[nf_arm_doce_top.scala 124:13]
  assign io_issue_sync = sync == 2'h2; // @[bfs_remote.scala 193:25]
  assign io_issue_sync_phase2 = sync == 2'h1; // @[bfs_remote.scala 194:32]
  assign io_remote_unvisited_size = unvisited_size_reg; // @[bfs_remote.scala 216:28]
  assign vertex_in_fifo_s_axis_aclk = clock; // @[bfs_remote.scala 183:48]
  assign vertex_in_fifo_s_axis_aresetn = ~reset; // @[bfs_remote.scala 184:39]
  assign vertex_in_fifo_s_axis_tdata = io_remote_in_w_bits_wdata; // @[bfs_remote.scala 187:34]
  assign vertex_in_fifo_s_axis_tkeep = io_remote_in_w_bits_wstrb; // @[bfs_remote.scala 186:34]
  assign vertex_in_fifo_s_axis_tlast = 1'h0;
  assign vertex_in_fifo_s_axis_tvalid = io_remote_in_w_valid; // @[bfs_remote.scala 185:35]
  assign vertex_in_fifo_s_axis_tid = 1'h0;
  assign vertex_in_fifo_m_axis_tready = is_sync | _vertex_in_fifo_io_m_axis_tready_T; // @[Mux.scala 98:16]
  always @(posedge clock) begin
    if (reset) begin // @[bfs_remote.scala 190:21]
      sync <= 2'h0; // @[bfs_remote.scala 190:21]
    end else if (is_sync) begin // @[bfs_remote.scala 195:16]
      sync <= _sync_T_1; // @[bfs_remote.scala 196:10]
    end else if (~io_start & io_signal) begin // @[bfs_remote.scala 197:37]
      sync <= 2'h0; // @[bfs_remote.scala 198:10]
    end
    if (reset) begin // @[bfs_remote.scala 210:35]
      unvisited_size_reg <= 32'h0; // @[bfs_remote.scala 210:35]
    end else if (is_sync) begin // @[bfs_remote.scala 211:16]
      unvisited_size_reg <= _unvisited_size_reg_T_2; // @[bfs_remote.scala 212:24]
    end else if (_T_1) begin // @[bfs_remote.scala 213:37]
      unvisited_size_reg <= 32'h0; // @[bfs_remote.scala 214:24]
    end
    if (reset) begin // @[bfs_remote.scala 221:28]
      packet_recv <= 32'h0; // @[bfs_remote.scala 221:28]
    end else if (io_remote_in_w_valid & io_remote_in_w_ready) begin // @[bfs_remote.scala 223:53]
      packet_recv <= _packet_recv_T_1; // @[bfs_remote.scala 224:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  unvisited_size_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  packet_recv = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BFS_ps(
  input          clock,
  input          reset,
  input  [63:0]  io_config_awaddr,
  input          io_config_awvalid,
  output         io_config_awready,
  input  [63:0]  io_config_araddr,
  input          io_config_arvalid,
  output         io_config_arready,
  input  [31:0]  io_config_wdata,
  input  [3:0]   io_config_wstrb,
  input          io_config_wvalid,
  output         io_config_wready,
  output [31:0]  io_config_rdata,
  output [1:0]   io_config_rresp,
  output         io_config_rvalid,
  input          io_config_rready,
  output [1:0]   io_config_bresp,
  output         io_config_bvalid,
  input          io_config_bready,
  input          io_PLmemory_0_aw_ready,
  output         io_PLmemory_0_aw_valid,
  output [63:0]  io_PLmemory_0_aw_bits_awaddr,
  output [6:0]   io_PLmemory_0_aw_bits_awid,
  output [7:0]   io_PLmemory_0_aw_bits_awlen,
  output [2:0]   io_PLmemory_0_aw_bits_awsize,
  output [1:0]   io_PLmemory_0_aw_bits_awburst,
  output         io_PLmemory_0_aw_bits_awlock,
  input          io_PLmemory_0_ar_ready,
  output         io_PLmemory_0_ar_valid,
  output [63:0]  io_PLmemory_0_ar_bits_araddr,
  output [6:0]   io_PLmemory_0_ar_bits_arid,
  output [7:0]   io_PLmemory_0_ar_bits_arlen,
  output [2:0]   io_PLmemory_0_ar_bits_arsize,
  output [1:0]   io_PLmemory_0_ar_bits_arburst,
  output         io_PLmemory_0_ar_bits_arlock,
  input          io_PLmemory_0_w_ready,
  output         io_PLmemory_0_w_valid,
  output [511:0] io_PLmemory_0_w_bits_wdata,
  output [63:0]  io_PLmemory_0_w_bits_wstrb,
  output         io_PLmemory_0_w_bits_wlast,
  output         io_PLmemory_0_r_ready,
  input          io_PLmemory_0_r_valid,
  input  [511:0] io_PLmemory_0_r_bits_rdata,
  input  [6:0]   io_PLmemory_0_r_bits_rid,
  input          io_PLmemory_0_r_bits_rlast,
  output         io_PLmemory_0_b_ready,
  input          io_PLmemory_0_b_valid,
  input  [1:0]   io_PLmemory_0_b_bits_bresp,
  input  [6:0]   io_PLmemory_0_b_bits_bid,
  input          io_PLmemory_1_aw_ready,
  output         io_PLmemory_1_aw_valid,
  output [63:0]  io_PLmemory_1_aw_bits_awaddr,
  output [6:0]   io_PLmemory_1_aw_bits_awid,
  output [7:0]   io_PLmemory_1_aw_bits_awlen,
  output [2:0]   io_PLmemory_1_aw_bits_awsize,
  output [1:0]   io_PLmemory_1_aw_bits_awburst,
  output         io_PLmemory_1_aw_bits_awlock,
  input          io_PLmemory_1_ar_ready,
  output         io_PLmemory_1_ar_valid,
  output [63:0]  io_PLmemory_1_ar_bits_araddr,
  output [6:0]   io_PLmemory_1_ar_bits_arid,
  output [7:0]   io_PLmemory_1_ar_bits_arlen,
  output [2:0]   io_PLmemory_1_ar_bits_arsize,
  output [1:0]   io_PLmemory_1_ar_bits_arburst,
  output         io_PLmemory_1_ar_bits_arlock,
  input          io_PLmemory_1_w_ready,
  output         io_PLmemory_1_w_valid,
  output [511:0] io_PLmemory_1_w_bits_wdata,
  output [63:0]  io_PLmemory_1_w_bits_wstrb,
  output         io_PLmemory_1_w_bits_wlast,
  output         io_PLmemory_1_r_ready,
  input          io_PLmemory_1_r_valid,
  input  [511:0] io_PLmemory_1_r_bits_rdata,
  input  [6:0]   io_PLmemory_1_r_bits_rid,
  input          io_PLmemory_1_r_bits_rlast,
  output         io_PLmemory_1_b_ready,
  input          io_PLmemory_1_b_valid,
  input  [1:0]   io_PLmemory_1_b_bits_bresp,
  input  [6:0]   io_PLmemory_1_b_bits_bid,
  input          io_PSmemory_0_aw_ready,
  output         io_PSmemory_0_aw_valid,
  output [63:0]  io_PSmemory_0_aw_bits_awaddr,
  output [5:0]   io_PSmemory_0_aw_bits_awid,
  output [7:0]   io_PSmemory_0_aw_bits_awlen,
  output [2:0]   io_PSmemory_0_aw_bits_awsize,
  output [1:0]   io_PSmemory_0_aw_bits_awburst,
  output         io_PSmemory_0_aw_bits_awlock,
  input          io_PSmemory_0_ar_ready,
  output         io_PSmemory_0_ar_valid,
  output [63:0]  io_PSmemory_0_ar_bits_araddr,
  output [5:0]   io_PSmemory_0_ar_bits_arid,
  output [7:0]   io_PSmemory_0_ar_bits_arlen,
  output [2:0]   io_PSmemory_0_ar_bits_arsize,
  output [1:0]   io_PSmemory_0_ar_bits_arburst,
  output         io_PSmemory_0_ar_bits_arlock,
  input          io_PSmemory_0_w_ready,
  output         io_PSmemory_0_w_valid,
  output [127:0] io_PSmemory_0_w_bits_wdata,
  output [15:0]  io_PSmemory_0_w_bits_wstrb,
  output         io_PSmemory_0_w_bits_wlast,
  output         io_PSmemory_0_r_ready,
  input          io_PSmemory_0_r_valid,
  input  [127:0] io_PSmemory_0_r_bits_rdata,
  input  [5:0]   io_PSmemory_0_r_bits_rid,
  input          io_PSmemory_0_r_bits_rlast,
  output         io_PSmemory_0_b_ready,
  input          io_PSmemory_0_b_valid,
  input  [1:0]   io_PSmemory_0_b_bits_bresp,
  input  [5:0]   io_PSmemory_0_b_bits_bid,
  input          io_PSmemory_1_aw_ready,
  output         io_PSmemory_1_aw_valid,
  output [63:0]  io_PSmemory_1_aw_bits_awaddr,
  output [5:0]   io_PSmemory_1_aw_bits_awid,
  output [7:0]   io_PSmemory_1_aw_bits_awlen,
  output [2:0]   io_PSmemory_1_aw_bits_awsize,
  output [1:0]   io_PSmemory_1_aw_bits_awburst,
  output         io_PSmemory_1_aw_bits_awlock,
  input          io_PSmemory_1_ar_ready,
  output         io_PSmemory_1_ar_valid,
  output [63:0]  io_PSmemory_1_ar_bits_araddr,
  output [5:0]   io_PSmemory_1_ar_bits_arid,
  output [7:0]   io_PSmemory_1_ar_bits_arlen,
  output [2:0]   io_PSmemory_1_ar_bits_arsize,
  output [1:0]   io_PSmemory_1_ar_bits_arburst,
  output         io_PSmemory_1_ar_bits_arlock,
  input          io_PSmemory_1_w_ready,
  output         io_PSmemory_1_w_valid,
  output [127:0] io_PSmemory_1_w_bits_wdata,
  output [15:0]  io_PSmemory_1_w_bits_wstrb,
  output         io_PSmemory_1_w_bits_wlast,
  output         io_PSmemory_1_r_ready,
  input          io_PSmemory_1_r_valid,
  input  [127:0] io_PSmemory_1_r_bits_rdata,
  input  [5:0]   io_PSmemory_1_r_bits_rid,
  input          io_PSmemory_1_r_bits_rlast,
  output         io_PSmemory_1_b_ready,
  input          io_PSmemory_1_b_valid,
  input  [1:0]   io_PSmemory_1_b_bits_bresp,
  input  [5:0]   io_PSmemory_1_b_bits_bid,
  input          io_PSmemory_2_aw_ready,
  output         io_PSmemory_2_aw_valid,
  output [63:0]  io_PSmemory_2_aw_bits_awaddr,
  output [5:0]   io_PSmemory_2_aw_bits_awid,
  output [7:0]   io_PSmemory_2_aw_bits_awlen,
  output [2:0]   io_PSmemory_2_aw_bits_awsize,
  output [1:0]   io_PSmemory_2_aw_bits_awburst,
  output         io_PSmemory_2_aw_bits_awlock,
  input          io_PSmemory_2_ar_ready,
  output         io_PSmemory_2_ar_valid,
  output [63:0]  io_PSmemory_2_ar_bits_araddr,
  output [5:0]   io_PSmemory_2_ar_bits_arid,
  output [7:0]   io_PSmemory_2_ar_bits_arlen,
  output [2:0]   io_PSmemory_2_ar_bits_arsize,
  output [1:0]   io_PSmemory_2_ar_bits_arburst,
  output         io_PSmemory_2_ar_bits_arlock,
  input          io_PSmemory_2_w_ready,
  output         io_PSmemory_2_w_valid,
  output [127:0] io_PSmemory_2_w_bits_wdata,
  output [15:0]  io_PSmemory_2_w_bits_wstrb,
  output         io_PSmemory_2_w_bits_wlast,
  output         io_PSmemory_2_r_ready,
  input          io_PSmemory_2_r_valid,
  input  [127:0] io_PSmemory_2_r_bits_rdata,
  input  [5:0]   io_PSmemory_2_r_bits_rid,
  input          io_PSmemory_2_r_bits_rlast,
  output         io_PSmemory_2_b_ready,
  input          io_PSmemory_2_b_valid,
  input  [1:0]   io_PSmemory_2_b_bits_bresp,
  input  [5:0]   io_PSmemory_2_b_bits_bid,
  input          io_PSmemory_3_aw_ready,
  output         io_PSmemory_3_aw_valid,
  output [63:0]  io_PSmemory_3_aw_bits_awaddr,
  output [5:0]   io_PSmemory_3_aw_bits_awid,
  output [7:0]   io_PSmemory_3_aw_bits_awlen,
  output [2:0]   io_PSmemory_3_aw_bits_awsize,
  output [1:0]   io_PSmemory_3_aw_bits_awburst,
  output         io_PSmemory_3_aw_bits_awlock,
  input          io_PSmemory_3_ar_ready,
  output         io_PSmemory_3_ar_valid,
  output [63:0]  io_PSmemory_3_ar_bits_araddr,
  output [5:0]   io_PSmemory_3_ar_bits_arid,
  output [7:0]   io_PSmemory_3_ar_bits_arlen,
  output [2:0]   io_PSmemory_3_ar_bits_arsize,
  output [1:0]   io_PSmemory_3_ar_bits_arburst,
  output         io_PSmemory_3_ar_bits_arlock,
  input          io_PSmemory_3_w_ready,
  output         io_PSmemory_3_w_valid,
  output [127:0] io_PSmemory_3_w_bits_wdata,
  output [15:0]  io_PSmemory_3_w_bits_wstrb,
  output         io_PSmemory_3_w_bits_wlast,
  output         io_PSmemory_3_r_ready,
  input          io_PSmemory_3_r_valid,
  input  [127:0] io_PSmemory_3_r_bits_rdata,
  input  [5:0]   io_PSmemory_3_r_bits_rid,
  input          io_PSmemory_3_r_bits_rlast,
  output         io_PSmemory_3_b_ready,
  input          io_PSmemory_3_b_valid,
  input  [1:0]   io_PSmemory_3_b_bits_bresp,
  input  [5:0]   io_PSmemory_3_b_bits_bid,
  input          io_Re_memory_out_aw_ready,
  output         io_Re_memory_out_aw_valid,
  output [63:0]  io_Re_memory_out_aw_bits_awaddr,
  output [5:0]   io_Re_memory_out_aw_bits_awid,
  output [7:0]   io_Re_memory_out_aw_bits_awlen,
  output [2:0]   io_Re_memory_out_aw_bits_awsize,
  output [1:0]   io_Re_memory_out_aw_bits_awburst,
  output         io_Re_memory_out_aw_bits_awlock,
  input          io_Re_memory_out_ar_ready,
  output         io_Re_memory_out_ar_valid,
  output [63:0]  io_Re_memory_out_ar_bits_araddr,
  output [5:0]   io_Re_memory_out_ar_bits_arid,
  output [7:0]   io_Re_memory_out_ar_bits_arlen,
  output [2:0]   io_Re_memory_out_ar_bits_arsize,
  output [1:0]   io_Re_memory_out_ar_bits_arburst,
  output         io_Re_memory_out_ar_bits_arlock,
  input          io_Re_memory_out_w_ready,
  output         io_Re_memory_out_w_valid,
  output [511:0] io_Re_memory_out_w_bits_wdata,
  output [63:0]  io_Re_memory_out_w_bits_wstrb,
  output         io_Re_memory_out_w_bits_wlast,
  output         io_Re_memory_out_r_ready,
  input          io_Re_memory_out_r_valid,
  input  [511:0] io_Re_memory_out_r_bits_rdata,
  input  [5:0]   io_Re_memory_out_r_bits_rid,
  input          io_Re_memory_out_r_bits_rlast,
  output         io_Re_memory_out_b_ready,
  input          io_Re_memory_out_b_valid,
  input  [1:0]   io_Re_memory_out_b_bits_bresp,
  input  [5:0]   io_Re_memory_out_b_bits_bid,
  output         io_Re_memory_in_aw_ready,
  input          io_Re_memory_in_aw_valid,
  input  [63:0]  io_Re_memory_in_aw_bits_awaddr,
  input  [9:0]   io_Re_memory_in_aw_bits_awid,
  input  [7:0]   io_Re_memory_in_aw_bits_awlen,
  input  [2:0]   io_Re_memory_in_aw_bits_awsize,
  input  [1:0]   io_Re_memory_in_aw_bits_awburst,
  input          io_Re_memory_in_aw_bits_awlock,
  output         io_Re_memory_in_ar_ready,
  input          io_Re_memory_in_ar_valid,
  input  [63:0]  io_Re_memory_in_ar_bits_araddr,
  input  [9:0]   io_Re_memory_in_ar_bits_arid,
  input  [7:0]   io_Re_memory_in_ar_bits_arlen,
  input  [2:0]   io_Re_memory_in_ar_bits_arsize,
  input  [1:0]   io_Re_memory_in_ar_bits_arburst,
  input          io_Re_memory_in_ar_bits_arlock,
  output         io_Re_memory_in_w_ready,
  input          io_Re_memory_in_w_valid,
  input  [511:0] io_Re_memory_in_w_bits_wdata,
  input  [63:0]  io_Re_memory_in_w_bits_wstrb,
  input          io_Re_memory_in_w_bits_wlast,
  input          io_Re_memory_in_r_ready,
  output         io_Re_memory_in_r_valid,
  output [511:0] io_Re_memory_in_r_bits_rdata,
  output [9:0]   io_Re_memory_in_r_bits_rid,
  output         io_Re_memory_in_r_bits_rlast,
  input          io_Re_memory_in_b_ready,
  output         io_Re_memory_in_b_valid,
  output [1:0]   io_Re_memory_in_b_bits_bresp,
  output [9:0]   io_Re_memory_in_b_bits_bid
);
  wire  controls_clock; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_reset; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_0; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_1; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_2; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_3; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_4; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_5; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_6; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_7; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_8; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_9; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_10; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_11; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_16; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_17; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_data_18; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_0; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_1; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_2; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_3; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_4; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_5; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_6; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_7; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_8; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_9; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_10; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_11; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_12; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_13; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_14; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_15; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_fin_16; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_signal; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_start; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_level; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_unvisited_size; // @[nf_arm_doce_top_main.scala 35:24]
  wire [63:0] controls_io_traveled_edges; // @[nf_arm_doce_top_main.scala 35:24]
  wire [63:0] controls_io_config_awaddr; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_awvalid; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_awready; // @[nf_arm_doce_top_main.scala 35:24]
  wire [63:0] controls_io_config_araddr; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_arvalid; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_arready; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_config_wdata; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_wvalid; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_wready; // @[nf_arm_doce_top_main.scala 35:24]
  wire [31:0] controls_io_config_rdata; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_rvalid; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_rready; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_bvalid; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_config_bready; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_flush_cache; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_flush_cache_end; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_signal_ack; // @[nf_arm_doce_top_main.scala 35:24]
  wire  controls_io_performance_0; // @[nf_arm_doce_top_main.scala 35:24]
  wire  MemController_clock; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_reset; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_out_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_out_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [511:0] MemController_io_cacheable_out_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire [15:0] MemController_io_cacheable_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_0_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_0_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_0_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_1_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_1_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_1_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_2_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_2_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_2_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_3_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_3_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_3_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_4_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_4_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_4_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_5_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_5_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_5_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_6_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_6_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_6_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_7_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_7_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_7_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_8_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_8_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_8_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_9_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_9_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_9_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_10_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_10_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_10_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_11_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_11_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_11_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_12_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_12_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_12_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_13_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_13_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_13_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_14_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_14_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_14_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_15_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_cacheable_in_15_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_cacheable_in_15_bits_tdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_non_cacheable_in_aw_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_non_cacheable_in_aw_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [63:0] MemController_io_non_cacheable_in_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 38:29]
  wire [6:0] MemController_io_non_cacheable_in_aw_bits_awid; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_non_cacheable_in_w_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_non_cacheable_in_w_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [511:0] MemController_io_non_cacheable_in_w_bits_wdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire [63:0] MemController_io_non_cacheable_in_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_0_aw_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_0_aw_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [63:0] MemController_io_ddr_out_0_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_0_ar_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_0_ar_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [63:0] MemController_io_ddr_out_0_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_0_w_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_0_w_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [511:0] MemController_io_ddr_out_0_w_bits_wdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_0_w_bits_wlast; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_0_r_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [511:0] MemController_io_ddr_out_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_1_aw_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_1_aw_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [63:0] MemController_io_ddr_out_1_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 38:29]
  wire [6:0] MemController_io_ddr_out_1_aw_bits_awid; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_1_w_ready; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_ddr_out_1_w_valid; // @[nf_arm_doce_top_main.scala 38:29]
  wire [511:0] MemController_io_ddr_out_1_w_bits_wdata; // @[nf_arm_doce_top_main.scala 38:29]
  wire [63:0] MemController_io_ddr_out_1_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 38:29]
  wire [63:0] MemController_io_tiers_base_addr_0; // @[nf_arm_doce_top_main.scala 38:29]
  wire [63:0] MemController_io_tiers_base_addr_1; // @[nf_arm_doce_top_main.scala 38:29]
  wire [31:0] MemController_io_unvisited_size; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_start; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_signal; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_end; // @[nf_arm_doce_top_main.scala 38:29]
  wire  MemController_io_signal_ack; // @[nf_arm_doce_top_main.scala 38:29]
  wire  Applys_0_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_0_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_0_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_0_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_0_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_0_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_0_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_0_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_0_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_0_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_1_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_1_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_1_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_1_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_1_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_1_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_1_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_1_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_1_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_1_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_2_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_2_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_2_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_2_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_2_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_2_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_2_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_2_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_2_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_2_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_3_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_3_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_3_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_3_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_3_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_3_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_3_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_3_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_3_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_3_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_4_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_4_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_4_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_4_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_4_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_4_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_4_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_4_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_4_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_4_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_4_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_5_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_5_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_5_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_5_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_5_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_5_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_5_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_5_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_5_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_5_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_5_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_6_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_6_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_6_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_6_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_6_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_6_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_6_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_6_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_6_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_6_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_6_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_7_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_7_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_7_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_7_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_7_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_7_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_7_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_7_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_7_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_7_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_7_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_8_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_8_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_8_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_8_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_8_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_8_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_8_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_8_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_8_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_8_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_8_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_9_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_9_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_9_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_9_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_9_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_9_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_9_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_9_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_9_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_9_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_9_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_10_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_10_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_10_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_10_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_10_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_10_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_10_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_10_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_10_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_10_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_10_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_11_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_11_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_11_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_11_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_11_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_11_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_11_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_11_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_11_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_11_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_11_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_12_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_12_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_12_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_12_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_12_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_12_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_12_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_12_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_12_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_12_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_12_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_13_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_13_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_13_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_13_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_13_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_13_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_13_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_13_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_13_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_13_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_13_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_14_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_14_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_14_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_14_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_14_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_14_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_14_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_14_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_14_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_14_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_14_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_15_clock; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_15_reset; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_15_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_15_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [1023:0] Applys_15_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_15_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_15_io_ddr_out_ready; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_15_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 40:16]
  wire [31:0] Applys_15_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_15_io_end; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Applys_15_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 40:16]
  wire  Gathers_clock; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_reset; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_ddr_in_ready; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_ddr_in_valid; // @[nf_arm_doce_top_main.scala 42:23]
  wire [511:0] Gathers_io_ddr_in_bits_tdata; // @[nf_arm_doce_top_main.scala 42:23]
  wire [15:0] Gathers_io_ddr_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_0_ready; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_0_valid; // @[nf_arm_doce_top_main.scala 42:23]
  wire [31:0] Gathers_io_gather_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_1_ready; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_1_valid; // @[nf_arm_doce_top_main.scala 42:23]
  wire [31:0] Gathers_io_gather_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_2_ready; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_2_valid; // @[nf_arm_doce_top_main.scala 42:23]
  wire [31:0] Gathers_io_gather_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_3_ready; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_3_valid; // @[nf_arm_doce_top_main.scala 42:23]
  wire [31:0] Gathers_io_gather_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_4_ready; // @[nf_arm_doce_top_main.scala 42:23]
  wire  Gathers_io_gather_out_4_valid; // @[nf_arm_doce_top_main.scala 42:23]
  wire [31:0] Gathers_io_gather_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 42:23]
  wire  LevelCache_clock; // @[nf_arm_doce_top_main.scala 43:26]
  wire  LevelCache_reset; // @[nf_arm_doce_top_main.scala 43:26]
  wire  LevelCache_io_ddr_aw_ready; // @[nf_arm_doce_top_main.scala 43:26]
  wire  LevelCache_io_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 43:26]
  wire [63:0] LevelCache_io_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 43:26]
  wire [6:0] LevelCache_io_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 43:26]
  wire  LevelCache_io_ddr_w_ready; // @[nf_arm_doce_top_main.scala 43:26]
  wire  LevelCache_io_ddr_w_valid; // @[nf_arm_doce_top_main.scala 43:26]
  wire [511:0] LevelCache_io_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 43:26]
  wire [63:0] LevelCache_io_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 43:26]
  wire  LevelCache_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 43:26]
  wire  LevelCache_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 43:26]
  wire [31:0] LevelCache_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 43:26]
  wire [31:0] LevelCache_io_level; // @[nf_arm_doce_top_main.scala 43:26]
  wire [63:0] LevelCache_io_level_base_addr; // @[nf_arm_doce_top_main.scala 43:26]
  wire  LevelCache_io_end; // @[nf_arm_doce_top_main.scala 43:26]
  wire  LevelCache_io_flush; // @[nf_arm_doce_top_main.scala 43:26]
  wire  Scatters_0_clock; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_reset; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_0_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 45:16]
  wire [5:0] Scatters_0_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [7:0] Scatters_0_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 45:16]
  wire [2:0] Scatters_0_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [127:0] Scatters_0_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire [5:0] Scatters_0_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [31:0] Scatters_0_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [127:0] Scatters_0_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire [3:0] Scatters_0_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_0_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_0_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_signal; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_0_io_traveled_edges; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_start; // @[nf_arm_doce_top_main.scala 45:16]
  wire [31:0] Scatters_0_io_root; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_0_io_issue_sync; // @[nf_arm_doce_top_main.scala 45:16]
  wire [4:0] Scatters_0_io_recv_sync; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_clock; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_reset; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_1_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 45:16]
  wire [5:0] Scatters_1_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [7:0] Scatters_1_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 45:16]
  wire [2:0] Scatters_1_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [127:0] Scatters_1_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire [5:0] Scatters_1_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [31:0] Scatters_1_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [127:0] Scatters_1_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire [3:0] Scatters_1_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_1_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_1_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_signal; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_1_io_traveled_edges; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_1_io_issue_sync; // @[nf_arm_doce_top_main.scala 45:16]
  wire [4:0] Scatters_1_io_recv_sync; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_clock; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_reset; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_2_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 45:16]
  wire [5:0] Scatters_2_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [7:0] Scatters_2_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 45:16]
  wire [2:0] Scatters_2_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [127:0] Scatters_2_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire [5:0] Scatters_2_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [31:0] Scatters_2_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [127:0] Scatters_2_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire [3:0] Scatters_2_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_2_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_2_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_signal; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_2_io_traveled_edges; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_2_io_issue_sync; // @[nf_arm_doce_top_main.scala 45:16]
  wire [4:0] Scatters_2_io_recv_sync; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_clock; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_reset; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_ddr_ar_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_3_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 45:16]
  wire [5:0] Scatters_3_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [7:0] Scatters_3_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 45:16]
  wire [2:0] Scatters_3_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_ddr_r_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [127:0] Scatters_3_io_ddr_r_bits_rdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire [5:0] Scatters_3_io_ddr_r_bits_rid; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_ddr_r_bits_rlast; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_gather_in_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [31:0] Scatters_3_io_gather_in_bits_tdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 45:16]
  wire [127:0] Scatters_3_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 45:16]
  wire [3:0] Scatters_3_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_3_io_embedding_base_addr; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_3_io_edge_base_addr; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_signal; // @[nf_arm_doce_top_main.scala 45:16]
  wire [63:0] Scatters_3_io_traveled_edges; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Scatters_3_io_issue_sync; // @[nf_arm_doce_top_main.scala 45:16]
  wire [4:0] Scatters_3_io_recv_sync; // @[nf_arm_doce_top_main.scala 45:16]
  wire  Broadcaster_clock; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_reset; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_ddr_in_0_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_ddr_in_0_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [127:0] Broadcaster_io_ddr_in_0_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [3:0] Broadcaster_io_ddr_in_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_ddr_in_1_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_ddr_in_1_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [127:0] Broadcaster_io_ddr_in_1_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [3:0] Broadcaster_io_ddr_in_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_ddr_in_2_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_ddr_in_2_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [127:0] Broadcaster_io_ddr_in_2_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [3:0] Broadcaster_io_ddr_in_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_ddr_in_3_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_ddr_in_3_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [127:0] Broadcaster_io_ddr_in_3_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [3:0] Broadcaster_io_ddr_in_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_0_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_0_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_1_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_1_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_2_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_2_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_3_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_3_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_4_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_4_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_4_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_5_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_5_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_5_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_5_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_6_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_6_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_6_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_6_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_7_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_7_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_7_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_7_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_8_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_8_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_8_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_8_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_9_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_9_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_9_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_9_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_10_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_10_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_10_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_10_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_11_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_11_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_11_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_11_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_12_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_12_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_12_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_12_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_13_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_13_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_13_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_13_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_14_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_14_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_14_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_14_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_15_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_pe_out_15_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [1023:0] Broadcaster_io_pe_out_15_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [31:0] Broadcaster_io_pe_out_15_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_remote_out_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [511:0] Broadcaster_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [15:0] Broadcaster_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_remote_in_ready; // @[nf_arm_doce_top_main.scala 48:27]
  wire  Broadcaster_io_remote_in_valid; // @[nf_arm_doce_top_main.scala 48:27]
  wire [511:0] Broadcaster_io_remote_in_bits_tdata; // @[nf_arm_doce_top_main.scala 48:27]
  wire [15:0] Broadcaster_io_remote_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 48:27]
  wire  ReApply_clock; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_reset; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_xbar_in_valid; // @[nf_arm_doce_top_main.scala 49:23]
  wire [511:0] ReApply_io_xbar_in_bits_tdata; // @[nf_arm_doce_top_main.scala 49:23]
  wire [15:0] ReApply_io_xbar_in_bits_tkeep; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_remote_out_aw_ready; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_remote_out_aw_valid; // @[nf_arm_doce_top_main.scala 49:23]
  wire [63:0] ReApply_io_remote_out_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 49:23]
  wire [5:0] ReApply_io_remote_out_aw_bits_awid; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_remote_out_w_ready; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_remote_out_w_valid; // @[nf_arm_doce_top_main.scala 49:23]
  wire [511:0] ReApply_io_remote_out_w_bits_wdata; // @[nf_arm_doce_top_main.scala 49:23]
  wire [63:0] ReApply_io_remote_out_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 49:23]
  wire [3:0] ReApply_io_recv_sync; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_recv_sync_phase2; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_signal; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_signal_ack; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_local_fpga_id; // @[nf_arm_doce_top_main.scala 49:23]
  wire [63:0] ReApply_io_level_base_addr; // @[nf_arm_doce_top_main.scala 49:23]
  wire [31:0] ReApply_io_local_unvisited_size; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReApply_io_end; // @[nf_arm_doce_top_main.scala 49:23]
  wire  ReScatter_clock; // @[nf_arm_doce_top_main.scala 51:25]
  wire  ReScatter_reset; // @[nf_arm_doce_top_main.scala 51:25]
  wire  ReScatter_io_remote_in_w_ready; // @[nf_arm_doce_top_main.scala 51:25]
  wire  ReScatter_io_remote_in_w_valid; // @[nf_arm_doce_top_main.scala 51:25]
  wire [511:0] ReScatter_io_remote_in_w_bits_wdata; // @[nf_arm_doce_top_main.scala 51:25]
  wire [63:0] ReScatter_io_remote_in_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 51:25]
  wire  ReScatter_io_xbar_out_ready; // @[nf_arm_doce_top_main.scala 51:25]
  wire  ReScatter_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 51:25]
  wire [511:0] ReScatter_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 51:25]
  wire [15:0] ReScatter_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 51:25]
  wire  ReScatter_io_signal; // @[nf_arm_doce_top_main.scala 51:25]
  wire  ReScatter_io_start; // @[nf_arm_doce_top_main.scala 51:25]
  wire  ReScatter_io_issue_sync; // @[nf_arm_doce_top_main.scala 51:25]
  wire  ReScatter_io_issue_sync_phase2; // @[nf_arm_doce_top_main.scala 51:25]
  wire [31:0] ReScatter_io_remote_unvisited_size; // @[nf_arm_doce_top_main.scala 51:25]
  wire [63:0] _controls_io_traveled_edges_T_1 = Scatters_0_io_traveled_edges + Scatters_1_io_traveled_edges; // @[nf_arm_doce_top_main.scala 96:80]
  wire [63:0] _controls_io_traveled_edges_T_3 = _controls_io_traveled_edges_T_1 + Scatters_2_io_traveled_edges; // @[nf_arm_doce_top_main.scala 96:80]
  wire  _Scatters_0_io_recv_sync_WIRE_1 = Scatters_0_io_issue_sync; // @[nf_arm_doce_top_main.scala 117:32 nf_arm_doce_top_main.scala 117:32]
  wire  _Scatters_0_io_recv_sync_WIRE_0 = ReScatter_io_issue_sync; // @[nf_arm_doce_top_main.scala 117:32 nf_arm_doce_top_main.scala 117:32]
  wire [1:0] Scatters_0_io_recv_sync_lo = {_Scatters_0_io_recv_sync_WIRE_1,_Scatters_0_io_recv_sync_WIRE_0}; // @[nf_arm_doce_top_main.scala 117:103]
  wire  _Scatters_0_io_recv_sync_WIRE_4 = Scatters_3_io_issue_sync; // @[nf_arm_doce_top_main.scala 117:32 nf_arm_doce_top_main.scala 117:32]
  wire  _Scatters_0_io_recv_sync_WIRE_3 = Scatters_2_io_issue_sync; // @[nf_arm_doce_top_main.scala 117:32 nf_arm_doce_top_main.scala 117:32]
  wire [1:0] Scatters_0_io_recv_sync_hi_hi = {_Scatters_0_io_recv_sync_WIRE_4,_Scatters_0_io_recv_sync_WIRE_3}; // @[nf_arm_doce_top_main.scala 117:103]
  wire  _Scatters_0_io_recv_sync_WIRE_2 = Scatters_1_io_issue_sync; // @[nf_arm_doce_top_main.scala 117:32 nf_arm_doce_top_main.scala 117:32]
  wire [2:0] Scatters_0_io_recv_sync_hi = {_Scatters_0_io_recv_sync_WIRE_4,_Scatters_0_io_recv_sync_WIRE_3,
    _Scatters_0_io_recv_sync_WIRE_2}; // @[nf_arm_doce_top_main.scala 117:103]
  wire [1:0] ReApply_io_recv_sync_lo = {_Scatters_0_io_recv_sync_WIRE_2,_Scatters_0_io_recv_sync_WIRE_1}; // @[nf_arm_doce_top_main.scala 125:77]
  controller controls ( // @[nf_arm_doce_top_main.scala 35:24]
    .clock(controls_clock),
    .reset(controls_reset),
    .io_data_0(controls_io_data_0),
    .io_data_1(controls_io_data_1),
    .io_data_2(controls_io_data_2),
    .io_data_3(controls_io_data_3),
    .io_data_4(controls_io_data_4),
    .io_data_5(controls_io_data_5),
    .io_data_6(controls_io_data_6),
    .io_data_7(controls_io_data_7),
    .io_data_8(controls_io_data_8),
    .io_data_9(controls_io_data_9),
    .io_data_10(controls_io_data_10),
    .io_data_11(controls_io_data_11),
    .io_data_16(controls_io_data_16),
    .io_data_17(controls_io_data_17),
    .io_data_18(controls_io_data_18),
    .io_fin_0(controls_io_fin_0),
    .io_fin_1(controls_io_fin_1),
    .io_fin_2(controls_io_fin_2),
    .io_fin_3(controls_io_fin_3),
    .io_fin_4(controls_io_fin_4),
    .io_fin_5(controls_io_fin_5),
    .io_fin_6(controls_io_fin_6),
    .io_fin_7(controls_io_fin_7),
    .io_fin_8(controls_io_fin_8),
    .io_fin_9(controls_io_fin_9),
    .io_fin_10(controls_io_fin_10),
    .io_fin_11(controls_io_fin_11),
    .io_fin_12(controls_io_fin_12),
    .io_fin_13(controls_io_fin_13),
    .io_fin_14(controls_io_fin_14),
    .io_fin_15(controls_io_fin_15),
    .io_fin_16(controls_io_fin_16),
    .io_signal(controls_io_signal),
    .io_start(controls_io_start),
    .io_level(controls_io_level),
    .io_unvisited_size(controls_io_unvisited_size),
    .io_traveled_edges(controls_io_traveled_edges),
    .io_config_awaddr(controls_io_config_awaddr),
    .io_config_awvalid(controls_io_config_awvalid),
    .io_config_awready(controls_io_config_awready),
    .io_config_araddr(controls_io_config_araddr),
    .io_config_arvalid(controls_io_config_arvalid),
    .io_config_arready(controls_io_config_arready),
    .io_config_wdata(controls_io_config_wdata),
    .io_config_wvalid(controls_io_config_wvalid),
    .io_config_wready(controls_io_config_wready),
    .io_config_rdata(controls_io_config_rdata),
    .io_config_rvalid(controls_io_config_rvalid),
    .io_config_rready(controls_io_config_rready),
    .io_config_bvalid(controls_io_config_bvalid),
    .io_config_bready(controls_io_config_bready),
    .io_flush_cache(controls_io_flush_cache),
    .io_flush_cache_end(controls_io_flush_cache_end),
    .io_signal_ack(controls_io_signal_ack),
    .io_performance_0(controls_io_performance_0)
  );
  multi_port_mc MemController ( // @[nf_arm_doce_top_main.scala 38:29]
    .clock(MemController_clock),
    .reset(MemController_reset),
    .io_cacheable_out_ready(MemController_io_cacheable_out_ready),
    .io_cacheable_out_valid(MemController_io_cacheable_out_valid),
    .io_cacheable_out_bits_tdata(MemController_io_cacheable_out_bits_tdata),
    .io_cacheable_out_bits_tkeep(MemController_io_cacheable_out_bits_tkeep),
    .io_cacheable_in_0_ready(MemController_io_cacheable_in_0_ready),
    .io_cacheable_in_0_valid(MemController_io_cacheable_in_0_valid),
    .io_cacheable_in_0_bits_tdata(MemController_io_cacheable_in_0_bits_tdata),
    .io_cacheable_in_1_ready(MemController_io_cacheable_in_1_ready),
    .io_cacheable_in_1_valid(MemController_io_cacheable_in_1_valid),
    .io_cacheable_in_1_bits_tdata(MemController_io_cacheable_in_1_bits_tdata),
    .io_cacheable_in_2_ready(MemController_io_cacheable_in_2_ready),
    .io_cacheable_in_2_valid(MemController_io_cacheable_in_2_valid),
    .io_cacheable_in_2_bits_tdata(MemController_io_cacheable_in_2_bits_tdata),
    .io_cacheable_in_3_ready(MemController_io_cacheable_in_3_ready),
    .io_cacheable_in_3_valid(MemController_io_cacheable_in_3_valid),
    .io_cacheable_in_3_bits_tdata(MemController_io_cacheable_in_3_bits_tdata),
    .io_cacheable_in_4_ready(MemController_io_cacheable_in_4_ready),
    .io_cacheable_in_4_valid(MemController_io_cacheable_in_4_valid),
    .io_cacheable_in_4_bits_tdata(MemController_io_cacheable_in_4_bits_tdata),
    .io_cacheable_in_5_ready(MemController_io_cacheable_in_5_ready),
    .io_cacheable_in_5_valid(MemController_io_cacheable_in_5_valid),
    .io_cacheable_in_5_bits_tdata(MemController_io_cacheable_in_5_bits_tdata),
    .io_cacheable_in_6_ready(MemController_io_cacheable_in_6_ready),
    .io_cacheable_in_6_valid(MemController_io_cacheable_in_6_valid),
    .io_cacheable_in_6_bits_tdata(MemController_io_cacheable_in_6_bits_tdata),
    .io_cacheable_in_7_ready(MemController_io_cacheable_in_7_ready),
    .io_cacheable_in_7_valid(MemController_io_cacheable_in_7_valid),
    .io_cacheable_in_7_bits_tdata(MemController_io_cacheable_in_7_bits_tdata),
    .io_cacheable_in_8_ready(MemController_io_cacheable_in_8_ready),
    .io_cacheable_in_8_valid(MemController_io_cacheable_in_8_valid),
    .io_cacheable_in_8_bits_tdata(MemController_io_cacheable_in_8_bits_tdata),
    .io_cacheable_in_9_ready(MemController_io_cacheable_in_9_ready),
    .io_cacheable_in_9_valid(MemController_io_cacheable_in_9_valid),
    .io_cacheable_in_9_bits_tdata(MemController_io_cacheable_in_9_bits_tdata),
    .io_cacheable_in_10_ready(MemController_io_cacheable_in_10_ready),
    .io_cacheable_in_10_valid(MemController_io_cacheable_in_10_valid),
    .io_cacheable_in_10_bits_tdata(MemController_io_cacheable_in_10_bits_tdata),
    .io_cacheable_in_11_ready(MemController_io_cacheable_in_11_ready),
    .io_cacheable_in_11_valid(MemController_io_cacheable_in_11_valid),
    .io_cacheable_in_11_bits_tdata(MemController_io_cacheable_in_11_bits_tdata),
    .io_cacheable_in_12_ready(MemController_io_cacheable_in_12_ready),
    .io_cacheable_in_12_valid(MemController_io_cacheable_in_12_valid),
    .io_cacheable_in_12_bits_tdata(MemController_io_cacheable_in_12_bits_tdata),
    .io_cacheable_in_13_ready(MemController_io_cacheable_in_13_ready),
    .io_cacheable_in_13_valid(MemController_io_cacheable_in_13_valid),
    .io_cacheable_in_13_bits_tdata(MemController_io_cacheable_in_13_bits_tdata),
    .io_cacheable_in_14_ready(MemController_io_cacheable_in_14_ready),
    .io_cacheable_in_14_valid(MemController_io_cacheable_in_14_valid),
    .io_cacheable_in_14_bits_tdata(MemController_io_cacheable_in_14_bits_tdata),
    .io_cacheable_in_15_ready(MemController_io_cacheable_in_15_ready),
    .io_cacheable_in_15_valid(MemController_io_cacheable_in_15_valid),
    .io_cacheable_in_15_bits_tdata(MemController_io_cacheable_in_15_bits_tdata),
    .io_non_cacheable_in_aw_ready(MemController_io_non_cacheable_in_aw_ready),
    .io_non_cacheable_in_aw_valid(MemController_io_non_cacheable_in_aw_valid),
    .io_non_cacheable_in_aw_bits_awaddr(MemController_io_non_cacheable_in_aw_bits_awaddr),
    .io_non_cacheable_in_aw_bits_awid(MemController_io_non_cacheable_in_aw_bits_awid),
    .io_non_cacheable_in_w_ready(MemController_io_non_cacheable_in_w_ready),
    .io_non_cacheable_in_w_valid(MemController_io_non_cacheable_in_w_valid),
    .io_non_cacheable_in_w_bits_wdata(MemController_io_non_cacheable_in_w_bits_wdata),
    .io_non_cacheable_in_w_bits_wstrb(MemController_io_non_cacheable_in_w_bits_wstrb),
    .io_ddr_out_0_aw_ready(MemController_io_ddr_out_0_aw_ready),
    .io_ddr_out_0_aw_valid(MemController_io_ddr_out_0_aw_valid),
    .io_ddr_out_0_aw_bits_awaddr(MemController_io_ddr_out_0_aw_bits_awaddr),
    .io_ddr_out_0_ar_ready(MemController_io_ddr_out_0_ar_ready),
    .io_ddr_out_0_ar_valid(MemController_io_ddr_out_0_ar_valid),
    .io_ddr_out_0_ar_bits_araddr(MemController_io_ddr_out_0_ar_bits_araddr),
    .io_ddr_out_0_w_ready(MemController_io_ddr_out_0_w_ready),
    .io_ddr_out_0_w_valid(MemController_io_ddr_out_0_w_valid),
    .io_ddr_out_0_w_bits_wdata(MemController_io_ddr_out_0_w_bits_wdata),
    .io_ddr_out_0_w_bits_wlast(MemController_io_ddr_out_0_w_bits_wlast),
    .io_ddr_out_0_r_valid(MemController_io_ddr_out_0_r_valid),
    .io_ddr_out_0_r_bits_rdata(MemController_io_ddr_out_0_r_bits_rdata),
    .io_ddr_out_0_r_bits_rlast(MemController_io_ddr_out_0_r_bits_rlast),
    .io_ddr_out_1_aw_ready(MemController_io_ddr_out_1_aw_ready),
    .io_ddr_out_1_aw_valid(MemController_io_ddr_out_1_aw_valid),
    .io_ddr_out_1_aw_bits_awaddr(MemController_io_ddr_out_1_aw_bits_awaddr),
    .io_ddr_out_1_aw_bits_awid(MemController_io_ddr_out_1_aw_bits_awid),
    .io_ddr_out_1_w_ready(MemController_io_ddr_out_1_w_ready),
    .io_ddr_out_1_w_valid(MemController_io_ddr_out_1_w_valid),
    .io_ddr_out_1_w_bits_wdata(MemController_io_ddr_out_1_w_bits_wdata),
    .io_ddr_out_1_w_bits_wstrb(MemController_io_ddr_out_1_w_bits_wstrb),
    .io_tiers_base_addr_0(MemController_io_tiers_base_addr_0),
    .io_tiers_base_addr_1(MemController_io_tiers_base_addr_1),
    .io_unvisited_size(MemController_io_unvisited_size),
    .io_start(MemController_io_start),
    .io_signal(MemController_io_signal),
    .io_end(MemController_io_end),
    .io_signal_ack(MemController_io_signal_ack)
  );
  Scatter Applys_0 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_0_clock),
    .reset(Applys_0_reset),
    .io_xbar_in_ready(Applys_0_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_0_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_0_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_0_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_0_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_0_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_0_io_ddr_out_bits_tdata),
    .io_end(Applys_0_io_end),
    .io_local_fpga_id(Applys_0_io_local_fpga_id)
  );
  Scatter_1 Applys_1 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_1_clock),
    .reset(Applys_1_reset),
    .io_xbar_in_ready(Applys_1_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_1_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_1_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_1_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_1_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_1_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_1_io_ddr_out_bits_tdata),
    .io_end(Applys_1_io_end),
    .io_local_fpga_id(Applys_1_io_local_fpga_id)
  );
  Scatter_2 Applys_2 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_2_clock),
    .reset(Applys_2_reset),
    .io_xbar_in_ready(Applys_2_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_2_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_2_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_2_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_2_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_2_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_2_io_ddr_out_bits_tdata),
    .io_end(Applys_2_io_end),
    .io_local_fpga_id(Applys_2_io_local_fpga_id)
  );
  Scatter_3 Applys_3 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_3_clock),
    .reset(Applys_3_reset),
    .io_xbar_in_ready(Applys_3_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_3_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_3_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_3_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_3_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_3_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_3_io_ddr_out_bits_tdata),
    .io_end(Applys_3_io_end),
    .io_local_fpga_id(Applys_3_io_local_fpga_id)
  );
  Scatter_4 Applys_4 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_4_clock),
    .reset(Applys_4_reset),
    .io_xbar_in_ready(Applys_4_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_4_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_4_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_4_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_4_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_4_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_4_io_ddr_out_bits_tdata),
    .io_end(Applys_4_io_end),
    .io_local_fpga_id(Applys_4_io_local_fpga_id)
  );
  Scatter_5 Applys_5 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_5_clock),
    .reset(Applys_5_reset),
    .io_xbar_in_ready(Applys_5_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_5_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_5_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_5_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_5_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_5_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_5_io_ddr_out_bits_tdata),
    .io_end(Applys_5_io_end),
    .io_local_fpga_id(Applys_5_io_local_fpga_id)
  );
  Scatter_6 Applys_6 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_6_clock),
    .reset(Applys_6_reset),
    .io_xbar_in_ready(Applys_6_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_6_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_6_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_6_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_6_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_6_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_6_io_ddr_out_bits_tdata),
    .io_end(Applys_6_io_end),
    .io_local_fpga_id(Applys_6_io_local_fpga_id)
  );
  Scatter_7 Applys_7 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_7_clock),
    .reset(Applys_7_reset),
    .io_xbar_in_ready(Applys_7_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_7_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_7_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_7_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_7_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_7_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_7_io_ddr_out_bits_tdata),
    .io_end(Applys_7_io_end),
    .io_local_fpga_id(Applys_7_io_local_fpga_id)
  );
  Scatter_8 Applys_8 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_8_clock),
    .reset(Applys_8_reset),
    .io_xbar_in_ready(Applys_8_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_8_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_8_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_8_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_8_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_8_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_8_io_ddr_out_bits_tdata),
    .io_end(Applys_8_io_end),
    .io_local_fpga_id(Applys_8_io_local_fpga_id)
  );
  Scatter_9 Applys_9 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_9_clock),
    .reset(Applys_9_reset),
    .io_xbar_in_ready(Applys_9_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_9_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_9_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_9_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_9_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_9_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_9_io_ddr_out_bits_tdata),
    .io_end(Applys_9_io_end),
    .io_local_fpga_id(Applys_9_io_local_fpga_id)
  );
  Scatter_10 Applys_10 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_10_clock),
    .reset(Applys_10_reset),
    .io_xbar_in_ready(Applys_10_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_10_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_10_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_10_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_10_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_10_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_10_io_ddr_out_bits_tdata),
    .io_end(Applys_10_io_end),
    .io_local_fpga_id(Applys_10_io_local_fpga_id)
  );
  Scatter_11 Applys_11 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_11_clock),
    .reset(Applys_11_reset),
    .io_xbar_in_ready(Applys_11_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_11_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_11_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_11_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_11_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_11_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_11_io_ddr_out_bits_tdata),
    .io_end(Applys_11_io_end),
    .io_local_fpga_id(Applys_11_io_local_fpga_id)
  );
  Scatter_12 Applys_12 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_12_clock),
    .reset(Applys_12_reset),
    .io_xbar_in_ready(Applys_12_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_12_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_12_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_12_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_12_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_12_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_12_io_ddr_out_bits_tdata),
    .io_end(Applys_12_io_end),
    .io_local_fpga_id(Applys_12_io_local_fpga_id)
  );
  Scatter_13 Applys_13 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_13_clock),
    .reset(Applys_13_reset),
    .io_xbar_in_ready(Applys_13_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_13_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_13_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_13_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_13_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_13_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_13_io_ddr_out_bits_tdata),
    .io_end(Applys_13_io_end),
    .io_local_fpga_id(Applys_13_io_local_fpga_id)
  );
  Scatter_14 Applys_14 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_14_clock),
    .reset(Applys_14_reset),
    .io_xbar_in_ready(Applys_14_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_14_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_14_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_14_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_14_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_14_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_14_io_ddr_out_bits_tdata),
    .io_end(Applys_14_io_end),
    .io_local_fpga_id(Applys_14_io_local_fpga_id)
  );
  Scatter_15 Applys_15 ( // @[nf_arm_doce_top_main.scala 40:16]
    .clock(Applys_15_clock),
    .reset(Applys_15_reset),
    .io_xbar_in_ready(Applys_15_io_xbar_in_ready),
    .io_xbar_in_valid(Applys_15_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(Applys_15_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(Applys_15_io_xbar_in_bits_tkeep),
    .io_ddr_out_ready(Applys_15_io_ddr_out_ready),
    .io_ddr_out_valid(Applys_15_io_ddr_out_valid),
    .io_ddr_out_bits_tdata(Applys_15_io_ddr_out_bits_tdata),
    .io_end(Applys_15_io_end),
    .io_local_fpga_id(Applys_15_io_local_fpga_id)
  );
  Gather Gathers ( // @[nf_arm_doce_top_main.scala 42:23]
    .clock(Gathers_clock),
    .reset(Gathers_reset),
    .io_ddr_in_ready(Gathers_io_ddr_in_ready),
    .io_ddr_in_valid(Gathers_io_ddr_in_valid),
    .io_ddr_in_bits_tdata(Gathers_io_ddr_in_bits_tdata),
    .io_ddr_in_bits_tkeep(Gathers_io_ddr_in_bits_tkeep),
    .io_gather_out_0_ready(Gathers_io_gather_out_0_ready),
    .io_gather_out_0_valid(Gathers_io_gather_out_0_valid),
    .io_gather_out_0_bits_tdata(Gathers_io_gather_out_0_bits_tdata),
    .io_gather_out_1_ready(Gathers_io_gather_out_1_ready),
    .io_gather_out_1_valid(Gathers_io_gather_out_1_valid),
    .io_gather_out_1_bits_tdata(Gathers_io_gather_out_1_bits_tdata),
    .io_gather_out_2_ready(Gathers_io_gather_out_2_ready),
    .io_gather_out_2_valid(Gathers_io_gather_out_2_valid),
    .io_gather_out_2_bits_tdata(Gathers_io_gather_out_2_bits_tdata),
    .io_gather_out_3_ready(Gathers_io_gather_out_3_ready),
    .io_gather_out_3_valid(Gathers_io_gather_out_3_valid),
    .io_gather_out_3_bits_tdata(Gathers_io_gather_out_3_bits_tdata),
    .io_gather_out_4_ready(Gathers_io_gather_out_4_ready),
    .io_gather_out_4_valid(Gathers_io_gather_out_4_valid),
    .io_gather_out_4_bits_tdata(Gathers_io_gather_out_4_bits_tdata)
  );
  Apply LevelCache ( // @[nf_arm_doce_top_main.scala 43:26]
    .clock(LevelCache_clock),
    .reset(LevelCache_reset),
    .io_ddr_aw_ready(LevelCache_io_ddr_aw_ready),
    .io_ddr_aw_valid(LevelCache_io_ddr_aw_valid),
    .io_ddr_aw_bits_awaddr(LevelCache_io_ddr_aw_bits_awaddr),
    .io_ddr_aw_bits_awid(LevelCache_io_ddr_aw_bits_awid),
    .io_ddr_w_ready(LevelCache_io_ddr_w_ready),
    .io_ddr_w_valid(LevelCache_io_ddr_w_valid),
    .io_ddr_w_bits_wdata(LevelCache_io_ddr_w_bits_wdata),
    .io_ddr_w_bits_wstrb(LevelCache_io_ddr_w_bits_wstrb),
    .io_gather_in_ready(LevelCache_io_gather_in_ready),
    .io_gather_in_valid(LevelCache_io_gather_in_valid),
    .io_gather_in_bits_tdata(LevelCache_io_gather_in_bits_tdata),
    .io_level(LevelCache_io_level),
    .io_level_base_addr(LevelCache_io_level_base_addr),
    .io_end(LevelCache_io_end),
    .io_flush(LevelCache_io_flush)
  );
  Broadcast Scatters_0 ( // @[nf_arm_doce_top_main.scala 45:16]
    .clock(Scatters_0_clock),
    .reset(Scatters_0_reset),
    .io_ddr_ar_ready(Scatters_0_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_0_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_0_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_0_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_0_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_0_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_0_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_0_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_0_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_0_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_0_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_0_io_gather_in_ready),
    .io_gather_in_valid(Scatters_0_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_0_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_0_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_0_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_0_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_0_io_xbar_out_bits_tkeep),
    .io_embedding_base_addr(Scatters_0_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_0_io_edge_base_addr),
    .io_signal(Scatters_0_io_signal),
    .io_traveled_edges(Scatters_0_io_traveled_edges),
    .io_start(Scatters_0_io_start),
    .io_root(Scatters_0_io_root),
    .io_issue_sync(Scatters_0_io_issue_sync),
    .io_recv_sync(Scatters_0_io_recv_sync)
  );
  Broadcast_1 Scatters_1 ( // @[nf_arm_doce_top_main.scala 45:16]
    .clock(Scatters_1_clock),
    .reset(Scatters_1_reset),
    .io_ddr_ar_ready(Scatters_1_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_1_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_1_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_1_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_1_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_1_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_1_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_1_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_1_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_1_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_1_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_1_io_gather_in_ready),
    .io_gather_in_valid(Scatters_1_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_1_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_1_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_1_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_1_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_1_io_xbar_out_bits_tkeep),
    .io_embedding_base_addr(Scatters_1_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_1_io_edge_base_addr),
    .io_signal(Scatters_1_io_signal),
    .io_traveled_edges(Scatters_1_io_traveled_edges),
    .io_issue_sync(Scatters_1_io_issue_sync),
    .io_recv_sync(Scatters_1_io_recv_sync)
  );
  Broadcast_2 Scatters_2 ( // @[nf_arm_doce_top_main.scala 45:16]
    .clock(Scatters_2_clock),
    .reset(Scatters_2_reset),
    .io_ddr_ar_ready(Scatters_2_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_2_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_2_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_2_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_2_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_2_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_2_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_2_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_2_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_2_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_2_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_2_io_gather_in_ready),
    .io_gather_in_valid(Scatters_2_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_2_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_2_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_2_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_2_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_2_io_xbar_out_bits_tkeep),
    .io_embedding_base_addr(Scatters_2_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_2_io_edge_base_addr),
    .io_signal(Scatters_2_io_signal),
    .io_traveled_edges(Scatters_2_io_traveled_edges),
    .io_issue_sync(Scatters_2_io_issue_sync),
    .io_recv_sync(Scatters_2_io_recv_sync)
  );
  Broadcast_3 Scatters_3 ( // @[nf_arm_doce_top_main.scala 45:16]
    .clock(Scatters_3_clock),
    .reset(Scatters_3_reset),
    .io_ddr_ar_ready(Scatters_3_io_ddr_ar_ready),
    .io_ddr_ar_valid(Scatters_3_io_ddr_ar_valid),
    .io_ddr_ar_bits_araddr(Scatters_3_io_ddr_ar_bits_araddr),
    .io_ddr_ar_bits_arid(Scatters_3_io_ddr_ar_bits_arid),
    .io_ddr_ar_bits_arlen(Scatters_3_io_ddr_ar_bits_arlen),
    .io_ddr_ar_bits_arsize(Scatters_3_io_ddr_ar_bits_arsize),
    .io_ddr_r_ready(Scatters_3_io_ddr_r_ready),
    .io_ddr_r_valid(Scatters_3_io_ddr_r_valid),
    .io_ddr_r_bits_rdata(Scatters_3_io_ddr_r_bits_rdata),
    .io_ddr_r_bits_rid(Scatters_3_io_ddr_r_bits_rid),
    .io_ddr_r_bits_rlast(Scatters_3_io_ddr_r_bits_rlast),
    .io_gather_in_ready(Scatters_3_io_gather_in_ready),
    .io_gather_in_valid(Scatters_3_io_gather_in_valid),
    .io_gather_in_bits_tdata(Scatters_3_io_gather_in_bits_tdata),
    .io_xbar_out_ready(Scatters_3_io_xbar_out_ready),
    .io_xbar_out_valid(Scatters_3_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(Scatters_3_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(Scatters_3_io_xbar_out_bits_tkeep),
    .io_embedding_base_addr(Scatters_3_io_embedding_base_addr),
    .io_edge_base_addr(Scatters_3_io_edge_base_addr),
    .io_signal(Scatters_3_io_signal),
    .io_traveled_edges(Scatters_3_io_traveled_edges),
    .io_issue_sync(Scatters_3_io_issue_sync),
    .io_recv_sync(Scatters_3_io_recv_sync)
  );
  Remote_xbar Broadcaster ( // @[nf_arm_doce_top_main.scala 48:27]
    .clock(Broadcaster_clock),
    .reset(Broadcaster_reset),
    .io_ddr_in_0_ready(Broadcaster_io_ddr_in_0_ready),
    .io_ddr_in_0_valid(Broadcaster_io_ddr_in_0_valid),
    .io_ddr_in_0_bits_tdata(Broadcaster_io_ddr_in_0_bits_tdata),
    .io_ddr_in_0_bits_tkeep(Broadcaster_io_ddr_in_0_bits_tkeep),
    .io_ddr_in_1_ready(Broadcaster_io_ddr_in_1_ready),
    .io_ddr_in_1_valid(Broadcaster_io_ddr_in_1_valid),
    .io_ddr_in_1_bits_tdata(Broadcaster_io_ddr_in_1_bits_tdata),
    .io_ddr_in_1_bits_tkeep(Broadcaster_io_ddr_in_1_bits_tkeep),
    .io_ddr_in_2_ready(Broadcaster_io_ddr_in_2_ready),
    .io_ddr_in_2_valid(Broadcaster_io_ddr_in_2_valid),
    .io_ddr_in_2_bits_tdata(Broadcaster_io_ddr_in_2_bits_tdata),
    .io_ddr_in_2_bits_tkeep(Broadcaster_io_ddr_in_2_bits_tkeep),
    .io_ddr_in_3_ready(Broadcaster_io_ddr_in_3_ready),
    .io_ddr_in_3_valid(Broadcaster_io_ddr_in_3_valid),
    .io_ddr_in_3_bits_tdata(Broadcaster_io_ddr_in_3_bits_tdata),
    .io_ddr_in_3_bits_tkeep(Broadcaster_io_ddr_in_3_bits_tkeep),
    .io_pe_out_0_ready(Broadcaster_io_pe_out_0_ready),
    .io_pe_out_0_valid(Broadcaster_io_pe_out_0_valid),
    .io_pe_out_0_bits_tdata(Broadcaster_io_pe_out_0_bits_tdata),
    .io_pe_out_0_bits_tkeep(Broadcaster_io_pe_out_0_bits_tkeep),
    .io_pe_out_1_ready(Broadcaster_io_pe_out_1_ready),
    .io_pe_out_1_valid(Broadcaster_io_pe_out_1_valid),
    .io_pe_out_1_bits_tdata(Broadcaster_io_pe_out_1_bits_tdata),
    .io_pe_out_1_bits_tkeep(Broadcaster_io_pe_out_1_bits_tkeep),
    .io_pe_out_2_ready(Broadcaster_io_pe_out_2_ready),
    .io_pe_out_2_valid(Broadcaster_io_pe_out_2_valid),
    .io_pe_out_2_bits_tdata(Broadcaster_io_pe_out_2_bits_tdata),
    .io_pe_out_2_bits_tkeep(Broadcaster_io_pe_out_2_bits_tkeep),
    .io_pe_out_3_ready(Broadcaster_io_pe_out_3_ready),
    .io_pe_out_3_valid(Broadcaster_io_pe_out_3_valid),
    .io_pe_out_3_bits_tdata(Broadcaster_io_pe_out_3_bits_tdata),
    .io_pe_out_3_bits_tkeep(Broadcaster_io_pe_out_3_bits_tkeep),
    .io_pe_out_4_ready(Broadcaster_io_pe_out_4_ready),
    .io_pe_out_4_valid(Broadcaster_io_pe_out_4_valid),
    .io_pe_out_4_bits_tdata(Broadcaster_io_pe_out_4_bits_tdata),
    .io_pe_out_4_bits_tkeep(Broadcaster_io_pe_out_4_bits_tkeep),
    .io_pe_out_5_ready(Broadcaster_io_pe_out_5_ready),
    .io_pe_out_5_valid(Broadcaster_io_pe_out_5_valid),
    .io_pe_out_5_bits_tdata(Broadcaster_io_pe_out_5_bits_tdata),
    .io_pe_out_5_bits_tkeep(Broadcaster_io_pe_out_5_bits_tkeep),
    .io_pe_out_6_ready(Broadcaster_io_pe_out_6_ready),
    .io_pe_out_6_valid(Broadcaster_io_pe_out_6_valid),
    .io_pe_out_6_bits_tdata(Broadcaster_io_pe_out_6_bits_tdata),
    .io_pe_out_6_bits_tkeep(Broadcaster_io_pe_out_6_bits_tkeep),
    .io_pe_out_7_ready(Broadcaster_io_pe_out_7_ready),
    .io_pe_out_7_valid(Broadcaster_io_pe_out_7_valid),
    .io_pe_out_7_bits_tdata(Broadcaster_io_pe_out_7_bits_tdata),
    .io_pe_out_7_bits_tkeep(Broadcaster_io_pe_out_7_bits_tkeep),
    .io_pe_out_8_ready(Broadcaster_io_pe_out_8_ready),
    .io_pe_out_8_valid(Broadcaster_io_pe_out_8_valid),
    .io_pe_out_8_bits_tdata(Broadcaster_io_pe_out_8_bits_tdata),
    .io_pe_out_8_bits_tkeep(Broadcaster_io_pe_out_8_bits_tkeep),
    .io_pe_out_9_ready(Broadcaster_io_pe_out_9_ready),
    .io_pe_out_9_valid(Broadcaster_io_pe_out_9_valid),
    .io_pe_out_9_bits_tdata(Broadcaster_io_pe_out_9_bits_tdata),
    .io_pe_out_9_bits_tkeep(Broadcaster_io_pe_out_9_bits_tkeep),
    .io_pe_out_10_ready(Broadcaster_io_pe_out_10_ready),
    .io_pe_out_10_valid(Broadcaster_io_pe_out_10_valid),
    .io_pe_out_10_bits_tdata(Broadcaster_io_pe_out_10_bits_tdata),
    .io_pe_out_10_bits_tkeep(Broadcaster_io_pe_out_10_bits_tkeep),
    .io_pe_out_11_ready(Broadcaster_io_pe_out_11_ready),
    .io_pe_out_11_valid(Broadcaster_io_pe_out_11_valid),
    .io_pe_out_11_bits_tdata(Broadcaster_io_pe_out_11_bits_tdata),
    .io_pe_out_11_bits_tkeep(Broadcaster_io_pe_out_11_bits_tkeep),
    .io_pe_out_12_ready(Broadcaster_io_pe_out_12_ready),
    .io_pe_out_12_valid(Broadcaster_io_pe_out_12_valid),
    .io_pe_out_12_bits_tdata(Broadcaster_io_pe_out_12_bits_tdata),
    .io_pe_out_12_bits_tkeep(Broadcaster_io_pe_out_12_bits_tkeep),
    .io_pe_out_13_ready(Broadcaster_io_pe_out_13_ready),
    .io_pe_out_13_valid(Broadcaster_io_pe_out_13_valid),
    .io_pe_out_13_bits_tdata(Broadcaster_io_pe_out_13_bits_tdata),
    .io_pe_out_13_bits_tkeep(Broadcaster_io_pe_out_13_bits_tkeep),
    .io_pe_out_14_ready(Broadcaster_io_pe_out_14_ready),
    .io_pe_out_14_valid(Broadcaster_io_pe_out_14_valid),
    .io_pe_out_14_bits_tdata(Broadcaster_io_pe_out_14_bits_tdata),
    .io_pe_out_14_bits_tkeep(Broadcaster_io_pe_out_14_bits_tkeep),
    .io_pe_out_15_ready(Broadcaster_io_pe_out_15_ready),
    .io_pe_out_15_valid(Broadcaster_io_pe_out_15_valid),
    .io_pe_out_15_bits_tdata(Broadcaster_io_pe_out_15_bits_tdata),
    .io_pe_out_15_bits_tkeep(Broadcaster_io_pe_out_15_bits_tkeep),
    .io_remote_out_ready(Broadcaster_io_remote_out_ready),
    .io_remote_out_valid(Broadcaster_io_remote_out_valid),
    .io_remote_out_bits_tdata(Broadcaster_io_remote_out_bits_tdata),
    .io_remote_out_bits_tkeep(Broadcaster_io_remote_out_bits_tkeep),
    .io_remote_in_ready(Broadcaster_io_remote_in_ready),
    .io_remote_in_valid(Broadcaster_io_remote_in_valid),
    .io_remote_in_bits_tdata(Broadcaster_io_remote_in_bits_tdata),
    .io_remote_in_bits_tkeep(Broadcaster_io_remote_in_bits_tkeep)
  );
  Remote_Apply ReApply ( // @[nf_arm_doce_top_main.scala 49:23]
    .clock(ReApply_clock),
    .reset(ReApply_reset),
    .io_xbar_in_ready(ReApply_io_xbar_in_ready),
    .io_xbar_in_valid(ReApply_io_xbar_in_valid),
    .io_xbar_in_bits_tdata(ReApply_io_xbar_in_bits_tdata),
    .io_xbar_in_bits_tkeep(ReApply_io_xbar_in_bits_tkeep),
    .io_remote_out_aw_ready(ReApply_io_remote_out_aw_ready),
    .io_remote_out_aw_valid(ReApply_io_remote_out_aw_valid),
    .io_remote_out_aw_bits_awaddr(ReApply_io_remote_out_aw_bits_awaddr),
    .io_remote_out_aw_bits_awid(ReApply_io_remote_out_aw_bits_awid),
    .io_remote_out_w_ready(ReApply_io_remote_out_w_ready),
    .io_remote_out_w_valid(ReApply_io_remote_out_w_valid),
    .io_remote_out_w_bits_wdata(ReApply_io_remote_out_w_bits_wdata),
    .io_remote_out_w_bits_wstrb(ReApply_io_remote_out_w_bits_wstrb),
    .io_recv_sync(ReApply_io_recv_sync),
    .io_recv_sync_phase2(ReApply_io_recv_sync_phase2),
    .io_signal(ReApply_io_signal),
    .io_signal_ack(ReApply_io_signal_ack),
    .io_local_fpga_id(ReApply_io_local_fpga_id),
    .io_level_base_addr(ReApply_io_level_base_addr),
    .io_local_unvisited_size(ReApply_io_local_unvisited_size),
    .io_end(ReApply_io_end)
  );
  Remote_Scatter ReScatter ( // @[nf_arm_doce_top_main.scala 51:25]
    .clock(ReScatter_clock),
    .reset(ReScatter_reset),
    .io_remote_in_w_ready(ReScatter_io_remote_in_w_ready),
    .io_remote_in_w_valid(ReScatter_io_remote_in_w_valid),
    .io_remote_in_w_bits_wdata(ReScatter_io_remote_in_w_bits_wdata),
    .io_remote_in_w_bits_wstrb(ReScatter_io_remote_in_w_bits_wstrb),
    .io_xbar_out_ready(ReScatter_io_xbar_out_ready),
    .io_xbar_out_valid(ReScatter_io_xbar_out_valid),
    .io_xbar_out_bits_tdata(ReScatter_io_xbar_out_bits_tdata),
    .io_xbar_out_bits_tkeep(ReScatter_io_xbar_out_bits_tkeep),
    .io_signal(ReScatter_io_signal),
    .io_start(ReScatter_io_start),
    .io_issue_sync(ReScatter_io_issue_sync),
    .io_issue_sync_phase2(ReScatter_io_issue_sync_phase2),
    .io_remote_unvisited_size(ReScatter_io_remote_unvisited_size)
  );
  assign io_config_awready = controls_io_config_awready; // @[nf_arm_doce_top_main.scala 95:22]
  assign io_config_arready = controls_io_config_arready; // @[nf_arm_doce_top_main.scala 95:22]
  assign io_config_wready = controls_io_config_wready; // @[nf_arm_doce_top_main.scala 95:22]
  assign io_config_rdata = controls_io_config_rdata; // @[nf_arm_doce_top_main.scala 95:22]
  assign io_config_rresp = 2'h0; // @[nf_arm_doce_top_main.scala 95:22]
  assign io_config_rvalid = controls_io_config_rvalid; // @[nf_arm_doce_top_main.scala 95:22]
  assign io_config_bresp = 2'h0; // @[nf_arm_doce_top_main.scala 95:22]
  assign io_config_bvalid = controls_io_config_bvalid; // @[nf_arm_doce_top_main.scala 95:22]
  assign io_PLmemory_0_aw_valid = MemController_io_ddr_out_0_aw_valid; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_aw_bits_awaddr = MemController_io_ddr_out_0_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_aw_bits_awid = 7'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_aw_bits_awlen = 8'hf; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_aw_bits_awsize = 3'h6; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_ar_valid = MemController_io_ddr_out_0_ar_valid; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_ar_bits_araddr = MemController_io_ddr_out_0_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_ar_bits_arid = 7'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_ar_bits_arlen = 8'hf; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_ar_bits_arsize = 3'h6; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_w_valid = MemController_io_ddr_out_0_w_valid; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_w_bits_wdata = MemController_io_ddr_out_0_w_bits_wdata; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_w_bits_wstrb = 64'hffffffffffffffff; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_w_bits_wlast = MemController_io_ddr_out_0_w_bits_wlast; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_r_ready = 1'h1; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_0_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_aw_valid = MemController_io_ddr_out_1_aw_valid; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_aw_bits_awaddr = MemController_io_ddr_out_1_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_aw_bits_awid = MemController_io_ddr_out_1_aw_bits_awid; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_aw_bits_awsize = 3'h2; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_ar_valid = 1'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_ar_bits_araddr = 64'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_ar_bits_arid = 7'h40; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_ar_bits_arlen = 8'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_ar_bits_arsize = 3'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_ar_bits_arburst = 2'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_w_valid = MemController_io_ddr_out_1_w_valid; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_w_bits_wdata = MemController_io_ddr_out_1_w_bits_wdata; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_w_bits_wstrb = MemController_io_ddr_out_1_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_w_bits_wlast = 1'h1; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_r_ready = 1'h0; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PLmemory_1_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 54:15]
  assign io_PSmemory_0_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 85:18]
  assign io_PSmemory_0_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 46:12]
  assign io_PSmemory_0_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 47:10]
  assign io_PSmemory_0_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 48:11]
  assign io_PSmemory_0_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 49:12]
  assign io_PSmemory_0_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 50:13]
  assign io_PSmemory_0_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_0_ar_valid = Scatters_0_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_0_ar_bits_araddr = Scatters_0_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_0_ar_bits_arid = Scatters_0_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_0_ar_bits_arlen = Scatters_0_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_0_ar_bits_arsize = Scatters_0_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_0_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_0_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_0_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 87:17]
  assign io_PSmemory_0_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 61:11]
  assign io_PSmemory_0_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 62:11]
  assign io_PSmemory_0_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 63:11]
  assign io_PSmemory_0_r_ready = Scatters_0_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 63:18]
  assign io_PSmemory_0_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 83:17]
  assign io_PSmemory_1_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 85:18]
  assign io_PSmemory_1_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 46:12]
  assign io_PSmemory_1_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 47:10]
  assign io_PSmemory_1_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 48:11]
  assign io_PSmemory_1_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 49:12]
  assign io_PSmemory_1_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 50:13]
  assign io_PSmemory_1_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_1_ar_valid = Scatters_1_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_1_ar_bits_araddr = Scatters_1_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_1_ar_bits_arid = Scatters_1_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_1_ar_bits_arlen = Scatters_1_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_1_ar_bits_arsize = Scatters_1_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_1_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_1_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_1_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 87:17]
  assign io_PSmemory_1_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 61:11]
  assign io_PSmemory_1_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 62:11]
  assign io_PSmemory_1_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 63:11]
  assign io_PSmemory_1_r_ready = Scatters_1_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 63:18]
  assign io_PSmemory_1_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 83:17]
  assign io_PSmemory_2_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 85:18]
  assign io_PSmemory_2_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 46:12]
  assign io_PSmemory_2_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 47:10]
  assign io_PSmemory_2_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 48:11]
  assign io_PSmemory_2_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 49:12]
  assign io_PSmemory_2_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 50:13]
  assign io_PSmemory_2_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_2_ar_valid = Scatters_2_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_2_ar_bits_araddr = Scatters_2_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_2_ar_bits_arid = Scatters_2_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_2_ar_bits_arlen = Scatters_2_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_2_ar_bits_arsize = Scatters_2_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_2_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_2_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_2_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 87:17]
  assign io_PSmemory_2_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 61:11]
  assign io_PSmemory_2_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 62:11]
  assign io_PSmemory_2_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 63:11]
  assign io_PSmemory_2_r_ready = Scatters_2_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 63:18]
  assign io_PSmemory_2_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 83:17]
  assign io_PSmemory_3_aw_valid = 1'h0; // @[nf_arm_doce_top_main.scala 85:18]
  assign io_PSmemory_3_aw_bits_awaddr = 64'h0; // @[nf_arm_doce_top.scala 46:12]
  assign io_PSmemory_3_aw_bits_awid = 6'h0; // @[nf_arm_doce_top.scala 47:10]
  assign io_PSmemory_3_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top.scala 48:11]
  assign io_PSmemory_3_aw_bits_awsize = 3'h0; // @[nf_arm_doce_top.scala 49:12]
  assign io_PSmemory_3_aw_bits_awburst = 2'h0; // @[nf_arm_doce_top.scala 50:13]
  assign io_PSmemory_3_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top.scala 51:12]
  assign io_PSmemory_3_ar_valid = Scatters_3_io_ddr_ar_valid; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_3_ar_bits_araddr = Scatters_3_io_ddr_ar_bits_araddr; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_3_ar_bits_arid = Scatters_3_io_ddr_ar_bits_arid; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_3_ar_bits_arlen = Scatters_3_io_ddr_ar_bits_arlen; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_3_ar_bits_arsize = Scatters_3_io_ddr_ar_bits_arsize; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_3_ar_bits_arburst = 2'h1; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_3_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 64:19]
  assign io_PSmemory_3_w_valid = 1'h0; // @[nf_arm_doce_top_main.scala 87:17]
  assign io_PSmemory_3_w_bits_wdata = 128'h0; // @[nf_arm_doce_top.scala 61:11]
  assign io_PSmemory_3_w_bits_wstrb = 16'h0; // @[nf_arm_doce_top.scala 62:11]
  assign io_PSmemory_3_w_bits_wlast = 1'h0; // @[nf_arm_doce_top.scala 63:11]
  assign io_PSmemory_3_r_ready = Scatters_3_io_ddr_r_ready; // @[nf_arm_doce_top_main.scala 63:18]
  assign io_PSmemory_3_b_ready = 1'h0; // @[nf_arm_doce_top_main.scala 83:17]
  assign io_Re_memory_out_aw_valid = ReApply_io_remote_out_aw_valid; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_aw_bits_awaddr = ReApply_io_remote_out_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_aw_bits_awid = ReApply_io_remote_out_aw_bits_awid; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_aw_bits_awlen = 8'h0; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_aw_bits_awsize = 3'h6; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_aw_bits_awburst = 2'h1; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_aw_bits_awlock = 1'h0; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_ar_valid = 1'h0; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_ar_bits_araddr = 64'h0; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_ar_bits_arid = 6'h0; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_ar_bits_arlen = 8'h0; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_ar_bits_arsize = 3'h0; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_ar_bits_arburst = 2'h0; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_ar_bits_arlock = 1'h0; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_w_valid = ReApply_io_remote_out_w_valid; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_w_bits_wdata = ReApply_io_remote_out_w_bits_wdata; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_w_bits_wstrb = ReApply_io_remote_out_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_w_bits_wlast = 1'h1; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_r_ready = 1'h1; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_out_b_ready = 1'h1; // @[nf_arm_doce_top_main.scala 78:20]
  assign io_Re_memory_in_aw_ready = 1'h1; // @[nf_arm_doce_top_main.scala 76:26]
  assign io_Re_memory_in_ar_ready = 1'h0; // @[nf_arm_doce_top_main.scala 76:26]
  assign io_Re_memory_in_w_ready = ReScatter_io_remote_in_w_ready; // @[nf_arm_doce_top_main.scala 76:26]
  assign io_Re_memory_in_r_valid = 1'h0; // @[nf_arm_doce_top_main.scala 76:26]
  assign io_Re_memory_in_r_bits_rdata = 512'h0; // @[nf_arm_doce_top_main.scala 76:26]
  assign io_Re_memory_in_r_bits_rid = 10'h0; // @[nf_arm_doce_top_main.scala 76:26]
  assign io_Re_memory_in_r_bits_rlast = 1'h0; // @[nf_arm_doce_top_main.scala 76:26]
  assign io_Re_memory_in_b_valid = 1'h0; // @[nf_arm_doce_top_main.scala 76:26]
  assign io_Re_memory_in_b_bits_bresp = 2'h0; // @[nf_arm_doce_top_main.scala 76:26]
  assign io_Re_memory_in_b_bits_bid = 10'h0; // @[nf_arm_doce_top_main.scala 76:26]
  assign controls_clock = clock;
  assign controls_reset = reset;
  assign controls_io_fin_0 = Applys_0_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_1 = Applys_1_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_2 = Applys_2_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_3 = Applys_3_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_4 = Applys_4_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_5 = Applys_5_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_6 = Applys_6_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_7 = Applys_7_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_8 = Applys_8_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_9 = Applys_9_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_10 = Applys_10_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_11 = Applys_11_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_12 = Applys_12_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_13 = Applys_13_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_14 = Applys_14_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_15 = Applys_15_io_end; // @[nf_arm_doce_top_main.scala 72:26]
  assign controls_io_fin_16 = ReApply_io_end; // @[nf_arm_doce_top_main.scala 100:24]
  assign controls_io_unvisited_size = MemController_io_unvisited_size + ReScatter_io_remote_unvisited_size; // @[nf_arm_doce_top_main.scala 97:65]
  assign controls_io_traveled_edges = _controls_io_traveled_edges_T_3 + Scatters_3_io_traveled_edges; // @[nf_arm_doce_top_main.scala 96:80]
  assign controls_io_config_awaddr = io_config_awaddr; // @[nf_arm_doce_top_main.scala 95:22]
  assign controls_io_config_awvalid = io_config_awvalid; // @[nf_arm_doce_top_main.scala 95:22]
  assign controls_io_config_araddr = io_config_araddr; // @[nf_arm_doce_top_main.scala 95:22]
  assign controls_io_config_arvalid = io_config_arvalid; // @[nf_arm_doce_top_main.scala 95:22]
  assign controls_io_config_wdata = io_config_wdata; // @[nf_arm_doce_top_main.scala 95:22]
  assign controls_io_config_wvalid = io_config_wvalid; // @[nf_arm_doce_top_main.scala 95:22]
  assign controls_io_config_rready = io_config_rready; // @[nf_arm_doce_top_main.scala 95:22]
  assign controls_io_config_bready = io_config_bready; // @[nf_arm_doce_top_main.scala 95:22]
  assign controls_io_flush_cache_end = LevelCache_io_end; // @[nf_arm_doce_top_main.scala 98:31]
  assign controls_io_signal_ack = MemController_io_signal_ack & ReApply_io_signal_ack; // @[nf_arm_doce_top_main.scala 99:57]
  assign controls_io_performance_0 = ~ReApply_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 101:33]
  assign MemController_clock = clock;
  assign MemController_reset = reset;
  assign MemController_io_cacheable_out_ready = Gathers_io_ddr_in_ready; // @[nf_arm_doce_top_main.scala 55:21]
  assign MemController_io_cacheable_in_0_valid = Applys_0_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_0_bits_tdata = Applys_0_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_1_valid = Applys_1_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_1_bits_tdata = Applys_1_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_2_valid = Applys_2_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_2_bits_tdata = Applys_2_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_3_valid = Applys_3_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_3_bits_tdata = Applys_3_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_4_valid = Applys_4_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_4_bits_tdata = Applys_4_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_5_valid = Applys_5_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_5_bits_tdata = Applys_5_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_6_valid = Applys_6_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_6_bits_tdata = Applys_6_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_7_valid = Applys_7_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_7_bits_tdata = Applys_7_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_8_valid = Applys_8_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_8_bits_tdata = Applys_8_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_9_valid = Applys_9_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_9_bits_tdata = Applys_9_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_10_valid = Applys_10_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_10_bits_tdata = Applys_10_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_11_valid = Applys_11_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_11_bits_tdata = Applys_11_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_12_valid = Applys_12_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_12_bits_tdata = Applys_12_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_13_valid = Applys_13_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_13_bits_tdata = Applys_13_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_14_valid = Applys_14_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_14_bits_tdata = Applys_14_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_15_valid = Applys_15_io_ddr_out_valid; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_cacheable_in_15_bits_tdata = Applys_15_io_ddr_out_bits_tdata; // @[nf_arm_doce_top_main.scala 71:21]
  assign MemController_io_non_cacheable_in_aw_valid = LevelCache_io_ddr_aw_valid; // @[nf_arm_doce_top_main.scala 58:24]
  assign MemController_io_non_cacheable_in_aw_bits_awaddr = LevelCache_io_ddr_aw_bits_awaddr; // @[nf_arm_doce_top_main.scala 58:24]
  assign MemController_io_non_cacheable_in_aw_bits_awid = LevelCache_io_ddr_aw_bits_awid; // @[nf_arm_doce_top_main.scala 58:24]
  assign MemController_io_non_cacheable_in_w_valid = LevelCache_io_ddr_w_valid; // @[nf_arm_doce_top_main.scala 57:23]
  assign MemController_io_non_cacheable_in_w_bits_wdata = LevelCache_io_ddr_w_bits_wdata; // @[nf_arm_doce_top_main.scala 57:23]
  assign MemController_io_non_cacheable_in_w_bits_wstrb = LevelCache_io_ddr_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 57:23]
  assign MemController_io_ddr_out_0_aw_ready = io_PLmemory_0_aw_ready; // @[nf_arm_doce_top_main.scala 54:15]
  assign MemController_io_ddr_out_0_ar_ready = io_PLmemory_0_ar_ready; // @[nf_arm_doce_top_main.scala 54:15]
  assign MemController_io_ddr_out_0_w_ready = io_PLmemory_0_w_ready; // @[nf_arm_doce_top_main.scala 54:15]
  assign MemController_io_ddr_out_0_r_valid = io_PLmemory_0_r_valid; // @[nf_arm_doce_top_main.scala 54:15]
  assign MemController_io_ddr_out_0_r_bits_rdata = io_PLmemory_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 54:15]
  assign MemController_io_ddr_out_0_r_bits_rlast = io_PLmemory_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 54:15]
  assign MemController_io_ddr_out_1_aw_ready = io_PLmemory_1_aw_ready; // @[nf_arm_doce_top_main.scala 54:15]
  assign MemController_io_ddr_out_1_w_ready = io_PLmemory_1_w_ready; // @[nf_arm_doce_top_main.scala 54:15]
  assign MemController_io_tiers_base_addr_0 = {controls_io_data_9,controls_io_data_8}; // @[Cat.scala 30:58]
  assign MemController_io_tiers_base_addr_1 = {controls_io_data_11,controls_io_data_10}; // @[Cat.scala 30:58]
  assign MemController_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 123:26]
  assign MemController_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 122:27]
  assign MemController_io_end = controls_io_data_0[1]; // @[nf_arm_doce_top_main.scala 124:46]
  assign Applys_0_clock = clock;
  assign Applys_0_reset = reset;
  assign Applys_0_io_xbar_in_valid = Broadcaster_io_pe_out_0_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_0_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_0_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_0_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_0_io_ddr_out_ready = MemController_io_cacheable_in_0_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_0_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_1_clock = clock;
  assign Applys_1_reset = reset;
  assign Applys_1_io_xbar_in_valid = Broadcaster_io_pe_out_1_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_1_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_1_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_1_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_1_io_ddr_out_ready = MemController_io_cacheable_in_1_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_1_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_2_clock = clock;
  assign Applys_2_reset = reset;
  assign Applys_2_io_xbar_in_valid = Broadcaster_io_pe_out_2_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_2_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_2_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_2_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_2_io_ddr_out_ready = MemController_io_cacheable_in_2_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_2_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_3_clock = clock;
  assign Applys_3_reset = reset;
  assign Applys_3_io_xbar_in_valid = Broadcaster_io_pe_out_3_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_3_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_3_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_3_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_3_io_ddr_out_ready = MemController_io_cacheable_in_3_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_3_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_4_clock = clock;
  assign Applys_4_reset = reset;
  assign Applys_4_io_xbar_in_valid = Broadcaster_io_pe_out_4_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_4_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_4_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_4_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_4_io_ddr_out_ready = MemController_io_cacheable_in_4_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_4_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_5_clock = clock;
  assign Applys_5_reset = reset;
  assign Applys_5_io_xbar_in_valid = Broadcaster_io_pe_out_5_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_5_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_5_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_5_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_5_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_5_io_ddr_out_ready = MemController_io_cacheable_in_5_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_5_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_6_clock = clock;
  assign Applys_6_reset = reset;
  assign Applys_6_io_xbar_in_valid = Broadcaster_io_pe_out_6_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_6_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_6_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_6_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_6_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_6_io_ddr_out_ready = MemController_io_cacheable_in_6_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_6_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_7_clock = clock;
  assign Applys_7_reset = reset;
  assign Applys_7_io_xbar_in_valid = Broadcaster_io_pe_out_7_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_7_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_7_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_7_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_7_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_7_io_ddr_out_ready = MemController_io_cacheable_in_7_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_7_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_8_clock = clock;
  assign Applys_8_reset = reset;
  assign Applys_8_io_xbar_in_valid = Broadcaster_io_pe_out_8_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_8_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_8_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_8_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_8_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_8_io_ddr_out_ready = MemController_io_cacheable_in_8_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_8_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_9_clock = clock;
  assign Applys_9_reset = reset;
  assign Applys_9_io_xbar_in_valid = Broadcaster_io_pe_out_9_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_9_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_9_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_9_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_9_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_9_io_ddr_out_ready = MemController_io_cacheable_in_9_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_9_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_10_clock = clock;
  assign Applys_10_reset = reset;
  assign Applys_10_io_xbar_in_valid = Broadcaster_io_pe_out_10_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_10_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_10_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_10_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_10_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_10_io_ddr_out_ready = MemController_io_cacheable_in_10_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_10_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_11_clock = clock;
  assign Applys_11_reset = reset;
  assign Applys_11_io_xbar_in_valid = Broadcaster_io_pe_out_11_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_11_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_11_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_11_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_11_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_11_io_ddr_out_ready = MemController_io_cacheable_in_11_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_11_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_12_clock = clock;
  assign Applys_12_reset = reset;
  assign Applys_12_io_xbar_in_valid = Broadcaster_io_pe_out_12_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_12_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_12_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_12_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_12_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_12_io_ddr_out_ready = MemController_io_cacheable_in_12_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_12_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_13_clock = clock;
  assign Applys_13_reset = reset;
  assign Applys_13_io_xbar_in_valid = Broadcaster_io_pe_out_13_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_13_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_13_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_13_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_13_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_13_io_ddr_out_ready = MemController_io_cacheable_in_13_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_13_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_14_clock = clock;
  assign Applys_14_reset = reset;
  assign Applys_14_io_xbar_in_valid = Broadcaster_io_pe_out_14_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_14_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_14_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_14_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_14_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_14_io_ddr_out_ready = MemController_io_cacheable_in_14_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_14_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Applys_15_clock = clock;
  assign Applys_15_reset = reset;
  assign Applys_15_io_xbar_in_valid = Broadcaster_io_pe_out_15_valid; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_15_io_xbar_in_bits_tdata = Broadcaster_io_pe_out_15_bits_tdata; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_15_io_xbar_in_bits_tkeep = Broadcaster_io_pe_out_15_bits_tkeep; // @[nf_arm_doce_top_main.scala 70:21]
  assign Applys_15_io_ddr_out_ready = MemController_io_cacheable_in_15_ready; // @[nf_arm_doce_top_main.scala 71:21]
  assign Applys_15_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 131:38]
  assign Gathers_clock = clock;
  assign Gathers_reset = reset;
  assign Gathers_io_ddr_in_valid = MemController_io_cacheable_out_valid; // @[nf_arm_doce_top_main.scala 55:21]
  assign Gathers_io_ddr_in_bits_tdata = MemController_io_cacheable_out_bits_tdata; // @[nf_arm_doce_top_main.scala 55:21]
  assign Gathers_io_ddr_in_bits_tkeep = MemController_io_cacheable_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 55:21]
  assign Gathers_io_gather_out_0_ready = Scatters_0_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 62:22]
  assign Gathers_io_gather_out_1_ready = Scatters_1_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 62:22]
  assign Gathers_io_gather_out_2_ready = Scatters_2_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 62:22]
  assign Gathers_io_gather_out_3_ready = Scatters_3_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 62:22]
  assign Gathers_io_gather_out_4_ready = LevelCache_io_gather_in_ready; // @[nf_arm_doce_top_main.scala 56:27]
  assign LevelCache_clock = clock;
  assign LevelCache_reset = reset;
  assign LevelCache_io_ddr_aw_ready = MemController_io_non_cacheable_in_aw_ready; // @[nf_arm_doce_top_main.scala 58:24]
  assign LevelCache_io_ddr_w_ready = MemController_io_non_cacheable_in_w_ready; // @[nf_arm_doce_top_main.scala 57:23]
  assign LevelCache_io_gather_in_valid = Gathers_io_gather_out_4_valid; // @[nf_arm_doce_top_main.scala 56:27]
  assign LevelCache_io_gather_in_bits_tdata = Gathers_io_gather_out_4_bits_tdata; // @[nf_arm_doce_top_main.scala 56:27]
  assign LevelCache_io_level = controls_io_level; // @[nf_arm_doce_top_main.scala 105:23]
  assign LevelCache_io_level_base_addr = {controls_io_data_6,controls_io_data_5}; // @[Cat.scala 30:58]
  assign LevelCache_io_flush = controls_io_flush_cache; // @[nf_arm_doce_top_main.scala 103:23]
  assign Scatters_0_clock = clock;
  assign Scatters_0_reset = reset;
  assign Scatters_0_io_ddr_ar_ready = io_PSmemory_0_ar_ready; // @[nf_arm_doce_top_main.scala 64:19]
  assign Scatters_0_io_ddr_r_valid = io_PSmemory_0_r_valid; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_0_io_ddr_r_bits_rdata = io_PSmemory_0_r_bits_rdata; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_0_io_ddr_r_bits_rid = io_PSmemory_0_r_bits_rid; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_0_io_ddr_r_bits_rlast = io_PSmemory_0_r_bits_rlast; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_0_io_gather_in_valid = Gathers_io_gather_out_0_valid; // @[nf_arm_doce_top_main.scala 62:22]
  assign Scatters_0_io_gather_in_bits_tdata = Gathers_io_gather_out_0_bits_tdata; // @[nf_arm_doce_top_main.scala 62:22]
  assign Scatters_0_io_xbar_out_ready = Broadcaster_io_ddr_in_0_ready; // @[nf_arm_doce_top_main.scala 65:32]
  assign Scatters_0_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_0_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_0_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 109:19]
  assign Scatters_0_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 113:20]
  assign Scatters_0_io_root = controls_io_data_7; // @[nf_arm_doce_top_main.scala 108:17]
  assign Scatters_0_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 117:103]
  assign Scatters_1_clock = clock;
  assign Scatters_1_reset = reset;
  assign Scatters_1_io_ddr_ar_ready = io_PSmemory_1_ar_ready; // @[nf_arm_doce_top_main.scala 64:19]
  assign Scatters_1_io_ddr_r_valid = io_PSmemory_1_r_valid; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_1_io_ddr_r_bits_rdata = io_PSmemory_1_r_bits_rdata; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_1_io_ddr_r_bits_rid = io_PSmemory_1_r_bits_rid; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_1_io_ddr_r_bits_rlast = io_PSmemory_1_r_bits_rlast; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_1_io_gather_in_valid = Gathers_io_gather_out_1_valid; // @[nf_arm_doce_top_main.scala 62:22]
  assign Scatters_1_io_gather_in_bits_tdata = Gathers_io_gather_out_1_bits_tdata; // @[nf_arm_doce_top_main.scala 62:22]
  assign Scatters_1_io_xbar_out_ready = Broadcaster_io_ddr_in_1_ready; // @[nf_arm_doce_top_main.scala 65:32]
  assign Scatters_1_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_1_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_1_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 109:19]
  assign Scatters_1_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 117:103]
  assign Scatters_2_clock = clock;
  assign Scatters_2_reset = reset;
  assign Scatters_2_io_ddr_ar_ready = io_PSmemory_2_ar_ready; // @[nf_arm_doce_top_main.scala 64:19]
  assign Scatters_2_io_ddr_r_valid = io_PSmemory_2_r_valid; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_2_io_ddr_r_bits_rdata = io_PSmemory_2_r_bits_rdata; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_2_io_ddr_r_bits_rid = io_PSmemory_2_r_bits_rid; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_2_io_ddr_r_bits_rlast = io_PSmemory_2_r_bits_rlast; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_2_io_gather_in_valid = Gathers_io_gather_out_2_valid; // @[nf_arm_doce_top_main.scala 62:22]
  assign Scatters_2_io_gather_in_bits_tdata = Gathers_io_gather_out_2_bits_tdata; // @[nf_arm_doce_top_main.scala 62:22]
  assign Scatters_2_io_xbar_out_ready = Broadcaster_io_ddr_in_2_ready; // @[nf_arm_doce_top_main.scala 65:32]
  assign Scatters_2_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_2_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_2_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 109:19]
  assign Scatters_2_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 117:103]
  assign Scatters_3_clock = clock;
  assign Scatters_3_reset = reset;
  assign Scatters_3_io_ddr_ar_ready = io_PSmemory_3_ar_ready; // @[nf_arm_doce_top_main.scala 64:19]
  assign Scatters_3_io_ddr_r_valid = io_PSmemory_3_r_valid; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_3_io_ddr_r_bits_rdata = io_PSmemory_3_r_bits_rdata; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_3_io_ddr_r_bits_rid = io_PSmemory_3_r_bits_rid; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_3_io_ddr_r_bits_rlast = io_PSmemory_3_r_bits_rlast; // @[nf_arm_doce_top_main.scala 63:18]
  assign Scatters_3_io_gather_in_valid = Gathers_io_gather_out_3_valid; // @[nf_arm_doce_top_main.scala 62:22]
  assign Scatters_3_io_gather_in_bits_tdata = Gathers_io_gather_out_3_bits_tdata; // @[nf_arm_doce_top_main.scala 62:22]
  assign Scatters_3_io_xbar_out_ready = Broadcaster_io_ddr_in_3_ready; // @[nf_arm_doce_top_main.scala 65:32]
  assign Scatters_3_io_embedding_base_addr = {controls_io_data_2,controls_io_data_1}; // @[Cat.scala 30:58]
  assign Scatters_3_io_edge_base_addr = {controls_io_data_4,controls_io_data_3}; // @[Cat.scala 30:58]
  assign Scatters_3_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 109:19]
  assign Scatters_3_io_recv_sync = {Scatters_0_io_recv_sync_hi,Scatters_0_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 117:103]
  assign Broadcaster_clock = clock;
  assign Broadcaster_reset = reset;
  assign Broadcaster_io_ddr_in_0_valid = Scatters_0_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_0_bits_tdata = Scatters_0_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_0_bits_tkeep = Scatters_0_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_1_valid = Scatters_1_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_1_bits_tdata = Scatters_1_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_1_bits_tkeep = Scatters_1_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_2_valid = Scatters_2_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_2_bits_tdata = Scatters_2_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_2_bits_tkeep = Scatters_2_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_3_valid = Scatters_3_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_3_bits_tdata = Scatters_3_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_ddr_in_3_bits_tkeep = Scatters_3_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 65:32]
  assign Broadcaster_io_pe_out_0_ready = Applys_0_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_1_ready = Applys_1_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_2_ready = Applys_2_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_3_ready = Applys_3_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_4_ready = Applys_4_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_5_ready = Applys_5_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_6_ready = Applys_6_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_7_ready = Applys_7_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_8_ready = Applys_8_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_9_ready = Applys_9_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_10_ready = Applys_10_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_11_ready = Applys_11_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_12_ready = Applys_12_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_13_ready = Applys_13_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_14_ready = Applys_14_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_pe_out_15_ready = Applys_15_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 70:21]
  assign Broadcaster_io_remote_out_ready = ReApply_io_xbar_in_ready; // @[nf_arm_doce_top_main.scala 77:22]
  assign Broadcaster_io_remote_in_valid = ReScatter_io_xbar_out_valid; // @[nf_arm_doce_top_main.scala 75:28]
  assign Broadcaster_io_remote_in_bits_tdata = ReScatter_io_xbar_out_bits_tdata; // @[nf_arm_doce_top_main.scala 75:28]
  assign Broadcaster_io_remote_in_bits_tkeep = ReScatter_io_xbar_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 75:28]
  assign ReApply_clock = clock;
  assign ReApply_reset = reset;
  assign ReApply_io_xbar_in_valid = Broadcaster_io_remote_out_valid; // @[nf_arm_doce_top_main.scala 77:22]
  assign ReApply_io_xbar_in_bits_tdata = Broadcaster_io_remote_out_bits_tdata; // @[nf_arm_doce_top_main.scala 77:22]
  assign ReApply_io_xbar_in_bits_tkeep = Broadcaster_io_remote_out_bits_tkeep; // @[nf_arm_doce_top_main.scala 77:22]
  assign ReApply_io_remote_out_aw_ready = io_Re_memory_out_aw_ready; // @[nf_arm_doce_top_main.scala 78:20]
  assign ReApply_io_remote_out_w_ready = io_Re_memory_out_w_ready; // @[nf_arm_doce_top_main.scala 78:20]
  assign ReApply_io_recv_sync = {Scatters_0_io_recv_sync_hi_hi,ReApply_io_recv_sync_lo}; // @[nf_arm_doce_top_main.scala 125:77]
  assign ReApply_io_recv_sync_phase2 = ReScatter_io_issue_sync_phase2; // @[nf_arm_doce_top_main.scala 130:31]
  assign ReApply_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 128:21]
  assign ReApply_io_local_fpga_id = controls_io_data_16[0]; // @[nf_arm_doce_top_main.scala 126:28]
  assign ReApply_io_level_base_addr = {controls_io_data_18,controls_io_data_17}; // @[Cat.scala 30:58]
  assign ReApply_io_local_unvisited_size = MemController_io_unvisited_size; // @[nf_arm_doce_top_main.scala 129:35]
  assign ReScatter_clock = clock;
  assign ReScatter_reset = reset;
  assign ReScatter_io_remote_in_w_valid = io_Re_memory_in_w_valid; // @[nf_arm_doce_top_main.scala 76:26]
  assign ReScatter_io_remote_in_w_bits_wdata = io_Re_memory_in_w_bits_wdata; // @[nf_arm_doce_top_main.scala 76:26]
  assign ReScatter_io_remote_in_w_bits_wstrb = io_Re_memory_in_w_bits_wstrb; // @[nf_arm_doce_top_main.scala 76:26]
  assign ReScatter_io_xbar_out_ready = Broadcaster_io_remote_in_ready; // @[nf_arm_doce_top_main.scala 75:28]
  assign ReScatter_io_signal = controls_io_signal; // @[nf_arm_doce_top_main.scala 133:23]
  assign ReScatter_io_start = controls_io_start; // @[nf_arm_doce_top_main.scala 132:22]
endmodule
