`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/16/2022 09:57:13 AM
// Design Name: 
// Module Name: bfs_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bfs_top(
    input gt_txusrclk,
    input peripheral_reset,
    input doceclk,
    input cmacclk,
    
    input  [63:0]  io_config_awaddr,
  input          io_config_awvalid,
  output         io_config_awready,
  input  [63:0]  io_config_araddr,
  input          io_config_arvalid,
  output         io_config_arready,
  input  [31:0]  io_config_wdata,
  input  [3:0]   io_config_wstrb,
  input          io_config_wvalid,
  output         io_config_wready,
  output [31:0]  io_config_rdata,
  output [1:0]   io_config_rresp,
  output         io_config_rvalid,
  input          io_config_rready,
  output [1:0]   io_config_bresp,
  output         io_config_bvalid,
  input          io_config_bready,

  input [511:0]doce_axis_rxd_tdata,
  input [63:0]doce_axis_rxd_tkeep,
  input doce_axis_rxd_tlast,
  output doce_axis_rxd_tready,
  input doce_axis_rxd_tvalid,
  output [511:0]doce_axis_txd_tdata,
  output [63:0]doce_axis_txd_tkeep,
  output doce_axis_txd_tlast,
  input doce_axis_txd_tready,
  output doce_axis_txd_tvalid
    );

    wire [63:0]  io_PLmemory_awaddr;
    wire [5:0]   io_PLmemory_awid;
    wire [7:0]   io_PLmemory_awlen;
    wire [2:0]   io_PLmemory_awsize;
    wire [1:0]   io_PLmemory_awburst;
    wire         io_PLmemory_awlock;
    wire         io_PLmemory_awvalid;
    wire         io_PLmemory_awready;
    wire [63:0]  io_PLmemory_araddr;
    wire [5:0]   io_PLmemory_arid;
    wire [7:0]   io_PLmemory_arlen;
    wire [2:0]   io_PLmemory_arsize;
    wire [1:0]   io_PLmemory_arburst;
    wire         io_PLmemory_arlock;
    wire         io_PLmemory_arvalid;
    wire         io_PLmemory_arready;
    wire [511:0] io_PLmemory_wdata;
    wire [63:0]  io_PLmemory_wstrb;
    wire         io_PLmemory_wlast;
    wire         io_PLmemory_wvalid;
    wire         io_PLmemory_wready;
    wire  [511:0]io_PLmemory_rdata;
    wire  [5:0]  io_PLmemory_rid;
    wire         io_PLmemory_rlast;
    wire  [1:0]  io_PLmemory_rresp;
    wire         io_PLmemory_rvalid;
    wire         io_PLmemory_rready;
    wire  [1:0]  io_PLmemory_bresp;
    wire  [5:0]  io_PLmemory_bid;
    wire         io_PLmemory_bvalid;
    wire         io_PLmemory_bready;

    memory u_pl_memory(
    .gt_txusrclk(gt_txusrclk),
    .peripheral_reset(peripheral_reset),
    .M00_AXI_AWID           (io_PLmemory_awid),     
    .M00_AXI_AWADDR         (io_PLmemory_awaddr),   
    .M00_AXI_AWLEN          (io_PLmemory_awlen),    
    .M00_AXI_AWSIZE         (io_PLmemory_awsize),   
    .M00_AXI_AWBURST        (io_PLmemory_awburst),  
    .M00_AXI_AWLOCK         (io_PLmemory_awlock),   
    .M00_AXI_AWCACHE        (),  
    .M00_AXI_AWPROT         (),   
    .M00_AXI_AWVALID        (io_PLmemory_awvalid),  
    .M00_AXI_AWREADY        (io_PLmemory_awready), 
    .M00_AXI_WDATA          (io_PLmemory_wdata),    
    .M00_AXI_WSTRB          (io_PLmemory_wstrb),    
    .M00_AXI_WLAST          (io_PLmemory_wlast),    
    .M00_AXI_WVALID         (io_PLmemory_wvalid),   
    .M00_AXI_WREADY         (io_PLmemory_wready),  
    .M00_AXI_BID            (io_PLmemory_bid),     
    .M00_AXI_BRESP          (io_PLmemory_bresp),   
    .M00_AXI_BVALID         (io_PLmemory_bvalid),  
    .M00_AXI_BREADY         (io_PLmemory_bready),   
    .M00_AXI_ARID           (io_PLmemory_arid),     
    .M00_AXI_ARADDR         (io_PLmemory_araddr),   
    .M00_AXI_ARLEN          (io_PLmemory_arlen),    
    .M00_AXI_ARSIZE         (io_PLmemory_arsize),   
    .M00_AXI_ARBURST        (io_PLmemory_arburst),  
    .M00_AXI_ARLOCK         (io_PLmemory_arlock),   
    .M00_AXI_ARCACHE        (),  
    .M00_AXI_ARPROT         (),   
    .M00_AXI_ARVALID        (io_PLmemory_arvalid),  
    .M00_AXI_ARREADY        (io_PLmemory_arready), 
    .M00_AXI_RID            (io_PLmemory_rid),     
    .M00_AXI_RDATA          (io_PLmemory_rdata),   
    .M00_AXI_RRESP          (io_PLmemory_rresp),   
    .M00_AXI_RLAST          (io_PLmemory_rlast),   
    .M00_AXI_RVALID         (io_PLmemory_rvalid),  
    .M00_AXI_RREADY         (io_PLmemory_rready),   
                  
    .M01_AXI_AWID           (io_PLmemory_awid),        
    .M01_AXI_AWADDR         (io_PLmemory_awaddr),    
    .M01_AXI_AWLEN          (io_PLmemory_awlen),      
    .M01_AXI_AWSIZE         (io_PLmemory_awsize),    
    .M01_AXI_AWBURST        (io_PLmemory_awburst),  
    .M01_AXI_AWLOCK         (io_PLmemory_awlock),    
    .M01_AXI_AWCACHE        (),                       
    .M01_AXI_AWPROT         (),                        
    .M01_AXI_AWVALID        (io_PLmemory_awvalid),  
    .M01_AXI_AWREADY        (io_PLmemory_awready), 
    .M01_AXI_WDATA          (io_PLmemory_wdata),      
    .M01_AXI_WSTRB          (io_PLmemory_wstrb),      
    .M01_AXI_WLAST          (io_PLmemory_wlast),      
    .M01_AXI_WVALID         (io_PLmemory_wvalid),    
    .M01_AXI_WREADY         (io_PLmemory_wready),   
    .M01_AXI_BID            (io_PLmemory_bid),         
    .M01_AXI_BRESP          (io_PLmemory_bresp),     
    .M01_AXI_BVALID         (io_PLmemory_bvalid),   
    .M01_AXI_BREADY         (io_PLmemory_bready),    
    .M01_AXI_ARID           (io_PLmemory_arid),        
    .M01_AXI_ARADDR         (io_PLmemory_araddr),    
    .M01_AXI_ARLEN          (io_PLmemory_arlen),      
    .M01_AXI_ARSIZE         (io_PLmemory_arsize),    
    .M01_AXI_ARBURST        (io_PLmemory_arburst),  
    .M01_AXI_ARLOCK         (io_PLmemory_arlock),    
    .M01_AXI_ARCACHE        (),                       
    .M01_AXI_ARPROT         (),                        
    .M01_AXI_ARVALID        (io_PLmemory_arvalid),  
    .M01_AXI_ARREADY        (io_PLmemory_arready), 
    .M01_AXI_RID            (io_PLmemory_rid),         
    .M01_AXI_RDATA          (io_PLmemory_rdata),     
    .M01_AXI_RRESP          (io_PLmemory_rresp),     
    .M01_AXI_RLAST          (io_PLmemory_rlast),     
    .M01_AXI_RVALID         (io_PLmemory_rvalid),   
    .M01_AXI_RREADY         (io_PLmemory_rready)
    );
    
    wire [63:0]  io_PSmemory_0_0_awaddr;
    wire [5:0]   io_PSmemory_0_0_awid;
    wire [7:0]   io_PSmemory_0_0_awlen;
    wire [2:0]   io_PSmemory_0_0_awsize;
    wire [1:0]   io_PSmemory_0_0_awburst;
    wire         io_PSmemory_0_0_awlock;
    wire         io_PSmemory_0_0_awvalid;
    wire         io_PSmemory_0_0_awready;
    wire [63:0]  io_PSmemory_0_0_araddr;
    wire [5:0]   io_PSmemory_0_0_arid;
    wire [7:0]   io_PSmemory_0_0_arlen;
    wire [2:0]   io_PSmemory_0_0_arsize;
    wire [1:0]   io_PSmemory_0_0_arburst;
    wire         io_PSmemory_0_0_arlock;
    wire         io_PSmemory_0_0_arvalid;
    wire         io_PSmemory_0_0_arready;
    wire [511:0] io_PSmemory_0_0_wdata;
    wire [63:0]  io_PSmemory_0_0_wstrb;
    wire         io_PSmemory_0_0_wlast;
    wire         io_PSmemory_0_0_wvalid;
    wire         io_PSmemory_0_0_wready;
    wire  [511:0]io_PSmemory_0_0_rdata;
    wire  [5:0]  io_PSmemory_0_0_rid;
    wire         io_PSmemory_0_0_rlast;
    wire  [1:0]  io_PSmemory_0_0_rresp;
    wire         io_PSmemory_0_0_rvalid;
    wire         io_PSmemory_0_0_rready;
    wire  [1:0]  io_PSmemory_0_0_bresp;
    wire  [5:0]  io_PSmemory_0_0_bid;
    wire         io_PSmemory_0_0_bvalid;
    wire         io_PSmemory_0_0_bready;

    wire [63:0]  io_PSmemory_0_1_awaddr;
    wire [5:0]   io_PSmemory_0_1_awid;
    wire [7:0]   io_PSmemory_0_1_awlen;
    wire [2:0]   io_PSmemory_0_1_awsize;
    wire [1:0]   io_PSmemory_0_1_awburst;
    wire         io_PSmemory_0_1_awlock;
    wire         io_PSmemory_0_1_awvalid;
    wire         io_PSmemory_0_1_awready;
    wire [63:0]  io_PSmemory_0_1_araddr;
    wire [5:0]   io_PSmemory_0_1_arid;
    wire [7:0]   io_PSmemory_0_1_arlen;
    wire [2:0]   io_PSmemory_0_1_arsize;
    wire [1:0]   io_PSmemory_0_1_arburst;
    wire         io_PSmemory_0_1_arlock;
    wire         io_PSmemory_0_1_arvalid;
    wire         io_PSmemory_0_1_arready;
    wire [511:0] io_PSmemory_0_1_wdata;
    wire [63:0]  io_PSmemory_0_1_wstrb;
    wire         io_PSmemory_0_1_wlast;
    wire         io_PSmemory_0_1_wvalid;
    wire         io_PSmemory_0_1_wready;
    wire  [511:0]io_PSmemory_0_1_rdata;
    wire  [5:0]  io_PSmemory_0_1_rid;
    wire         io_PSmemory_0_1_rlast;
    wire  [1:0]  io_PSmemory_0_1_rresp;
    wire         io_PSmemory_0_1_rvalid;
    wire         io_PSmemory_0_1_rready;
    wire  [1:0]  io_PSmemory_0_1_bresp;
    wire  [5:0]  io_PSmemory_0_1_bid;
    wire         io_PSmemory_0_1_bvalid;
    wire         io_PSmemory_0_1_bready;

    memory u_hp0_memory(
    .gt_txusrclk(gt_txusrclk),
    .peripheral_reset(peripheral_reset),
    .M00_AXI_AWID           (io_PSmemory_0_0_awid),     
    .M00_AXI_AWADDR         (io_PSmemory_0_0_awaddr),   
    .M00_AXI_AWLEN          (io_PSmemory_0_0_awlen),    
    .M00_AXI_AWSIZE         (io_PSmemory_0_0_awsize),   
    .M00_AXI_AWBURST        (io_PSmemory_0_0_awburst),  
    .M00_AXI_AWLOCK         (io_PSmemory_0_0_awlock),   
    .M00_AXI_AWCACHE        (),  
    .M00_AXI_AWPROT         (),   
    .M00_AXI_AWVALID        (io_PSmemory_0_0_awvalid),  
    .M00_AXI_AWREADY        (io_PSmemory_0_0_awready), 
    .M00_AXI_WDATA          (io_PSmemory_0_0_wdata),    
    .M00_AXI_WSTRB          (io_PSmemory_0_0_wstrb),    
    .M00_AXI_WLAST          (io_PSmemory_0_0_wlast),    
    .M00_AXI_WVALID         (io_PSmemory_0_0_wvalid),   
    .M00_AXI_WREADY         (io_PSmemory_0_0_wready),  
    .M00_AXI_BID            (io_PSmemory_0_0_bid),     
    .M00_AXI_BRESP          (io_PSmemory_0_0_bresp),   
    .M00_AXI_BVALID         (io_PSmemory_0_0_bvalid),  
    .M00_AXI_BREADY         (io_PSmemory_0_0_bready),   
    .M00_AXI_ARID           (io_PSmemory_0_0_arid),     
    .M00_AXI_ARADDR         (io_PSmemory_0_0_araddr),   
    .M00_AXI_ARLEN          (io_PSmemory_0_0_arlen),    
    .M00_AXI_ARSIZE         (io_PSmemory_0_0_arsize),   
    .M00_AXI_ARBURST        (io_PSmemory_0_0_arburst),  
    .M00_AXI_ARLOCK         (io_PSmemory_0_0_arlock),   
    .M00_AXI_ARCACHE        (),  
    .M00_AXI_ARPROT         (),   
    .M00_AXI_ARVALID        (io_PSmemory_0_0_arvalid),  
    .M00_AXI_ARREADY        (io_PSmemory_0_0_arready), 
    .M00_AXI_RID            (io_PSmemory_0_0_rid),     
    .M00_AXI_RDATA          (io_PSmemory_0_0_rdata),   
    .M00_AXI_RRESP          (io_PSmemory_0_0_rresp),   
    .M00_AXI_RLAST          (io_PSmemory_0_0_rlast),   
    .M00_AXI_RVALID         (io_PSmemory_0_0_rvalid),  
    .M00_AXI_RREADY         (io_PSmemory_0_0_rready),   
                  
    .M01_AXI_AWID           (io_PSmemory_0_1_awid),        
    .M01_AXI_AWADDR         (io_PSmemory_0_1_awaddr),    
    .M01_AXI_AWLEN          (io_PSmemory_0_1_awlen),      
    .M01_AXI_AWSIZE         (io_PSmemory_0_1_awsize),    
    .M01_AXI_AWBURST        (io_PSmemory_0_1_awburst),  
    .M01_AXI_AWLOCK         (io_PSmemory_0_1_awlock),    
    .M01_AXI_AWCACHE        (),                       
    .M01_AXI_AWPROT         (),                        
    .M01_AXI_AWVALID        (io_PSmemory_0_1_awvalid),  
    .M01_AXI_AWREADY        (io_PSmemory_0_1_awready), 
    .M01_AXI_WDATA          (io_PSmemory_0_1_wdata),      
    .M01_AXI_WSTRB          (io_PSmemory_0_1_wstrb),      
    .M01_AXI_WLAST          (io_PSmemory_0_1_wlast),      
    .M01_AXI_WVALID         (io_PSmemory_0_1_wvalid),    
    .M01_AXI_WREADY         (io_PSmemory_0_1_wready),   
    .M01_AXI_BID            (io_PSmemory_0_1_bid),         
    .M01_AXI_BRESP          (io_PSmemory_0_1_bresp),     
    .M01_AXI_BVALID         (io_PSmemory_0_1_bvalid),   
    .M01_AXI_BREADY         (io_PSmemory_0_1_bready),    
    .M01_AXI_ARID           (io_PSmemory_0_1_arid),        
    .M01_AXI_ARADDR         (io_PSmemory_0_1_araddr),    
    .M01_AXI_ARLEN          (io_PSmemory_0_1_arlen),      
    .M01_AXI_ARSIZE         (io_PSmemory_0_1_arsize),    
    .M01_AXI_ARBURST        (io_PSmemory_0_1_arburst),  
    .M01_AXI_ARLOCK         (io_PSmemory_0_1_arlock),    
    .M01_AXI_ARCACHE        (),                       
    .M01_AXI_ARPROT         (),                        
    .M01_AXI_ARVALID        (io_PSmemory_0_1_arvalid),  
    .M01_AXI_ARREADY        (io_PSmemory_0_1_arready), 
    .M01_AXI_RID            (io_PSmemory_0_1_rid),         
    .M01_AXI_RDATA          (io_PSmemory_0_1_rdata),     
    .M01_AXI_RRESP          (io_PSmemory_0_1_rresp),     
    .M01_AXI_RLAST          (io_PSmemory_0_1_rlast),     
    .M01_AXI_RVALID         (io_PSmemory_0_1_rvalid),   
    .M01_AXI_RREADY         (io_PSmemory_0_1_rready) 
    );
    
    wire [63:0]  io_PSmemory_1_0_awaddr;
    wire [5:0]   io_PSmemory_1_0_awid;
    wire [7:0]   io_PSmemory_1_0_awlen;
    wire [2:0]   io_PSmemory_1_0_awsize;
    wire [1:0]   io_PSmemory_1_0_awburst;
    wire         io_PSmemory_1_0_awlock;
    wire         io_PSmemory_1_0_awvalid;
    wire         io_PSmemory_1_0_awready;
    wire [63:0]  io_PSmemory_1_0_araddr;
    wire [5:0]   io_PSmemory_1_0_arid;
    wire [7:0]   io_PSmemory_1_0_arlen;
    wire [2:0]   io_PSmemory_1_0_arsize;
    wire [1:0]   io_PSmemory_1_0_arburst;
    wire         io_PSmemory_1_0_arlock;
    wire         io_PSmemory_1_0_arvalid;
    wire         io_PSmemory_1_0_arready;
    wire [511:0] io_PSmemory_1_0_wdata;
    wire [63:0]  io_PSmemory_1_0_wstrb;
    wire         io_PSmemory_1_0_wlast;
    wire         io_PSmemory_1_0_wvalid;
    wire         io_PSmemory_1_0_wready;
    wire  [511:0]io_PSmemory_1_0_rdata;
    wire  [5:0]  io_PSmemory_1_0_rid;
    wire         io_PSmemory_1_0_rlast;
    wire  [1:0]  io_PSmemory_1_0_rresp;
    wire         io_PSmemory_1_0_rvalid;
    wire         io_PSmemory_1_0_rready;
    wire  [1:0]  io_PSmemory_1_0_bresp;
    wire  [5:0]  io_PSmemory_1_0_bid;
    wire         io_PSmemory_1_0_bvalid;
    wire         io_PSmemory_1_0_bready;

    wire [63:0]  io_PSmemory_1_1_awaddr;
    wire [5:0]   io_PSmemory_1_1_awid;
    wire [7:0]   io_PSmemory_1_1_awlen;
    wire [2:0]   io_PSmemory_1_1_awsize;
    wire [1:0]   io_PSmemory_1_1_awburst;
    wire         io_PSmemory_1_1_awlock;
    wire         io_PSmemory_1_1_awvalid;
    wire         io_PSmemory_1_1_awready;
    wire [63:0]  io_PSmemory_1_1_araddr;
    wire [5:0]   io_PSmemory_1_1_arid;
    wire [7:0]   io_PSmemory_1_1_arlen;
    wire [2:0]   io_PSmemory_1_1_arsize;
    wire [1:0]   io_PSmemory_1_1_arburst;
    wire         io_PSmemory_1_1_arlock;
    wire         io_PSmemory_1_1_arvalid;
    wire         io_PSmemory_1_1_arready;
    wire [511:0] io_PSmemory_1_1_wdata;
    wire [63:0]  io_PSmemory_1_1_wstrb;
    wire         io_PSmemory_1_1_wlast;
    wire         io_PSmemory_1_1_wvalid;
    wire         io_PSmemory_1_1_wready;
    wire  [511:0]io_PSmemory_1_1_rdata;
    wire  [5:0]  io_PSmemory_1_1_rid;
    wire         io_PSmemory_1_1_rlast;
    wire  [1:0]  io_PSmemory_1_1_rresp;
    wire         io_PSmemory_1_1_rvalid;
    wire         io_PSmemory_1_1_rready;
    wire  [1:0]  io_PSmemory_1_1_bresp;
    wire  [5:0]  io_PSmemory_1_1_bid;
    wire         io_PSmemory_1_1_bvalid;
    wire         io_PSmemory_1_1_bready;

    memory u_hp1_memory(
    .gt_txusrclk(gt_txusrclk),
    .peripheral_reset(peripheral_reset),
    .M00_AXI_AWID           (io_PSmemory_1_0_awid),     
    .M00_AXI_AWADDR         (io_PSmemory_1_0_awaddr),   
    .M00_AXI_AWLEN          (io_PSmemory_1_0_awlen),    
    .M00_AXI_AWSIZE         (io_PSmemory_1_0_awsize),   
    .M00_AXI_AWBURST        (io_PSmemory_1_0_awburst),  
    .M00_AXI_AWLOCK         (io_PSmemory_1_0_awlock),   
    .M00_AXI_AWCACHE        (),  
    .M00_AXI_AWPROT         (),   
    .M00_AXI_AWVALID        (io_PSmemory_1_0_awvalid),  
    .M00_AXI_AWREADY        (io_PSmemory_1_0_awready), 
    .M00_AXI_WDATA          (io_PSmemory_1_0_wdata),    
    .M00_AXI_WSTRB          (io_PSmemory_1_0_wstrb),    
    .M00_AXI_WLAST          (io_PSmemory_1_0_wlast),    
    .M00_AXI_WVALID         (io_PSmemory_1_0_wvalid),   
    .M00_AXI_WREADY         (io_PSmemory_1_0_wready),  
    .M00_AXI_BID            (io_PSmemory_1_0_bid),     
    .M00_AXI_BRESP          (io_PSmemory_1_0_bresp),   
    .M00_AXI_BVALID         (io_PSmemory_1_0_bvalid),  
    .M00_AXI_BREADY         (io_PSmemory_1_0_bready),   
    .M00_AXI_ARID           (io_PSmemory_1_0_arid),     
    .M00_AXI_ARADDR         (io_PSmemory_1_0_araddr),   
    .M00_AXI_ARLEN          (io_PSmemory_1_0_arlen),    
    .M00_AXI_ARSIZE         (io_PSmemory_1_0_arsize),   
    .M00_AXI_ARBURST        (io_PSmemory_1_0_arburst),  
    .M00_AXI_ARLOCK         (io_PSmemory_1_0_arlock),   
    .M00_AXI_ARCACHE        (),  
    .M00_AXI_ARPROT         (),   
    .M00_AXI_ARVALID        (io_PSmemory_1_0_arvalid),  
    .M00_AXI_ARREADY        (io_PSmemory_1_0_arready), 
    .M00_AXI_RID            (io_PSmemory_1_0_rid),     
    .M00_AXI_RDATA          (io_PSmemory_1_0_rdata),   
    .M00_AXI_RRESP          (io_PSmemory_1_0_rresp),   
    .M00_AXI_RLAST          (io_PSmemory_1_0_rlast),   
    .M00_AXI_RVALID         (io_PSmemory_1_0_rvalid),  
    .M00_AXI_RREADY         (io_PSmemory_1_0_rready),   
                  
    .M01_AXI_AWID           (io_PSmemory_1_1_awid),        
    .M01_AXI_AWADDR         (io_PSmemory_1_1_awaddr),    
    .M01_AXI_AWLEN          (io_PSmemory_1_1_awlen),      
    .M01_AXI_AWSIZE         (io_PSmemory_1_1_awsize),    
    .M01_AXI_AWBURST        (io_PSmemory_1_1_awburst),  
    .M01_AXI_AWLOCK         (io_PSmemory_1_1_awlock),    
    .M01_AXI_AWCACHE        (),                       
    .M01_AXI_AWPROT         (),                        
    .M01_AXI_AWVALID        (io_PSmemory_1_1_awvalid),  
    .M01_AXI_AWREADY        (io_PSmemory_1_1_awready), 
    .M01_AXI_WDATA          (io_PSmemory_1_1_wdata),      
    .M01_AXI_WSTRB          (io_PSmemory_1_1_wstrb),      
    .M01_AXI_WLAST          (io_PSmemory_1_1_wlast),      
    .M01_AXI_WVALID         (io_PSmemory_1_1_wvalid),    
    .M01_AXI_WREADY         (io_PSmemory_1_1_wready),   
    .M01_AXI_BID            (io_PSmemory_1_1_bid),         
    .M01_AXI_BRESP          (io_PSmemory_1_1_bresp),     
    .M01_AXI_BVALID         (io_PSmemory_1_1_bvalid),   
    .M01_AXI_BREADY         (io_PSmemory_1_1_bready),    
    .M01_AXI_ARID           (io_PSmemory_1_1_arid),        
    .M01_AXI_ARADDR         (io_PSmemory_1_1_araddr),    
    .M01_AXI_ARLEN          (io_PSmemory_1_1_arlen),      
    .M01_AXI_ARSIZE         (io_PSmemory_1_1_arsize),    
    .M01_AXI_ARBURST        (io_PSmemory_1_1_arburst),  
    .M01_AXI_ARLOCK         (io_PSmemory_1_1_arlock),    
    .M01_AXI_ARCACHE        (),                       
    .M01_AXI_ARPROT         (),                        
    .M01_AXI_ARVALID        (io_PSmemory_1_1_arvalid),  
    .M01_AXI_ARREADY        (io_PSmemory_1_1_arready), 
    .M01_AXI_RID            (io_PSmemory_1_1_rid),         
    .M01_AXI_RDATA          (io_PSmemory_1_1_rdata),     
    .M01_AXI_RRESP          (io_PSmemory_1_1_rresp),     
    .M01_AXI_RLAST          (io_PSmemory_1_1_rlast),     
    .M01_AXI_RVALID         (io_PSmemory_1_1_rvalid),   
    .M01_AXI_RREADY         (io_PSmemory_1_1_rready) 
    );
    
    wire [63:0]  io_PSmemory_2_0_awaddr;
    wire [5:0]   io_PSmemory_2_0_awid;
    wire [7:0]   io_PSmemory_2_0_awlen;
    wire [2:0]   io_PSmemory_2_0_awsize;
    wire [1:0]   io_PSmemory_2_0_awburst;
    wire         io_PSmemory_2_0_awlock;
    wire         io_PSmemory_2_0_awvalid;
    wire         io_PSmemory_2_0_awready;
    wire [63:0]  io_PSmemory_2_0_araddr;
    wire [5:0]   io_PSmemory_2_0_arid;
    wire [7:0]   io_PSmemory_2_0_arlen;
    wire [2:0]   io_PSmemory_2_0_arsize;
    wire [1:0]   io_PSmemory_2_0_arburst;
    wire         io_PSmemory_2_0_arlock;
    wire         io_PSmemory_2_0_arvalid;
    wire         io_PSmemory_2_0_arready;
    wire [511:0] io_PSmemory_2_0_wdata;
    wire [63:0]  io_PSmemory_2_0_wstrb;
    wire         io_PSmemory_2_0_wlast;
    wire         io_PSmemory_2_0_wvalid;
    wire         io_PSmemory_2_0_wready;
    wire  [511:0]io_PSmemory_2_0_rdata;
    wire  [5:0]  io_PSmemory_2_0_rid;
    wire         io_PSmemory_2_0_rlast;
    wire  [1:0]  io_PSmemory_2_0_rresp;
    wire         io_PSmemory_2_0_rvalid;
    wire         io_PSmemory_2_0_rready;
    wire  [1:0]  io_PSmemory_2_0_bresp;
    wire  [5:0]  io_PSmemory_2_0_bid;
    wire         io_PSmemory_2_0_bvalid;
    wire         io_PSmemory_2_0_bready;

    wire [63:0]  io_PSmemory_2_1_awaddr;
    wire [5:0]   io_PSmemory_2_1_awid;
    wire [7:0]   io_PSmemory_2_1_awlen;
    wire [2:0]   io_PSmemory_2_1_awsize;
    wire [1:0]   io_PSmemory_2_1_awburst;
    wire         io_PSmemory_2_1_awlock;
    wire         io_PSmemory_2_1_awvalid;
    wire         io_PSmemory_2_1_awready;
    wire [63:0]  io_PSmemory_2_1_araddr;
    wire [5:0]   io_PSmemory_2_1_arid;
    wire [7:0]   io_PSmemory_2_1_arlen;
    wire [2:0]   io_PSmemory_2_1_arsize;
    wire [1:0]   io_PSmemory_2_1_arburst;
    wire         io_PSmemory_2_1_arlock;
    wire         io_PSmemory_2_1_arvalid;
    wire         io_PSmemory_2_1_arready;
    wire [511:0] io_PSmemory_2_1_wdata;
    wire [63:0]  io_PSmemory_2_1_wstrb;
    wire         io_PSmemory_2_1_wlast;
    wire         io_PSmemory_2_1_wvalid;
    wire         io_PSmemory_2_1_wready;
    wire  [511:0]io_PSmemory_2_1_rdata;
    wire  [5:0]  io_PSmemory_2_1_rid;
    wire         io_PSmemory_2_1_rlast;
    wire  [1:0]  io_PSmemory_2_1_rresp;
    wire         io_PSmemory_2_1_rvalid;
    wire         io_PSmemory_2_1_rready;
    wire  [1:0]  io_PSmemory_2_1_bresp;
    wire  [5:0]  io_PSmemory_2_1_bid;
    wire         io_PSmemory_2_1_bvalid;
    wire         io_PSmemory_2_1_bready;

    memory u_hp2_memory(
    .gt_txusrclk(gt_txusrclk),
    .peripheral_reset(peripheral_reset),
    .M00_AXI_AWID           (io_PSmemory_2_0_awid),     
    .M00_AXI_AWADDR         (io_PSmemory_2_0_awaddr),   
    .M00_AXI_AWLEN          (io_PSmemory_2_0_awlen),    
    .M00_AXI_AWSIZE         (io_PSmemory_2_0_awsize),   
    .M00_AXI_AWBURST        (io_PSmemory_2_0_awburst),  
    .M00_AXI_AWLOCK         (io_PSmemory_2_0_awlock),   
    .M00_AXI_AWCACHE        (),  
    .M00_AXI_AWPROT         (),   
    .M00_AXI_AWVALID        (io_PSmemory_2_0_awvalid),  
    .M00_AXI_AWREADY        (io_PSmemory_2_0_awready), 
    .M00_AXI_WDATA          (io_PSmemory_2_0_wdata),    
    .M00_AXI_WSTRB          (io_PSmemory_2_0_wstrb),    
    .M00_AXI_WLAST          (io_PSmemory_2_0_wlast),    
    .M00_AXI_WVALID         (io_PSmemory_2_0_wvalid),   
    .M00_AXI_WREADY         (io_PSmemory_2_0_wready),  
    .M00_AXI_BID            (io_PSmemory_2_0_bid),     
    .M00_AXI_BRESP          (io_PSmemory_2_0_bresp),   
    .M00_AXI_BVALID         (io_PSmemory_2_0_bvalid),  
    .M00_AXI_BREADY         (io_PSmemory_2_0_bready),   
    .M00_AXI_ARID           (io_PSmemory_2_0_arid),     
    .M00_AXI_ARADDR         (io_PSmemory_2_0_araddr),   
    .M00_AXI_ARLEN          (io_PSmemory_2_0_arlen),    
    .M00_AXI_ARSIZE         (io_PSmemory_2_0_arsize),   
    .M00_AXI_ARBURST        (io_PSmemory_2_0_arburst),  
    .M00_AXI_ARLOCK         (io_PSmemory_2_0_arlock),   
    .M00_AXI_ARCACHE        (),  
    .M00_AXI_ARPROT         (),   
    .M00_AXI_ARVALID        (io_PSmemory_2_0_arvalid),  
    .M00_AXI_ARREADY        (io_PSmemory_2_0_arready), 
    .M00_AXI_RID            (io_PSmemory_2_0_rid),     
    .M00_AXI_RDATA          (io_PSmemory_2_0_rdata),   
    .M00_AXI_RRESP          (io_PSmemory_2_0_rresp),   
    .M00_AXI_RLAST          (io_PSmemory_2_0_rlast),   
    .M00_AXI_RVALID         (io_PSmemory_2_0_rvalid),  
    .M00_AXI_RREADY         (io_PSmemory_2_0_rready),   
                  
    .M01_AXI_AWID           (io_PSmemory_2_1_awid),        
    .M01_AXI_AWADDR         (io_PSmemory_2_1_awaddr),    
    .M01_AXI_AWLEN          (io_PSmemory_2_1_awlen),      
    .M01_AXI_AWSIZE         (io_PSmemory_2_1_awsize),    
    .M01_AXI_AWBURST        (io_PSmemory_2_1_awburst),  
    .M01_AXI_AWLOCK         (io_PSmemory_2_1_awlock),    
    .M01_AXI_AWCACHE        (),                       
    .M01_AXI_AWPROT         (),                        
    .M01_AXI_AWVALID        (io_PSmemory_2_1_awvalid),  
    .M01_AXI_AWREADY        (io_PSmemory_2_1_awready), 
    .M01_AXI_WDATA          (io_PSmemory_2_1_wdata),      
    .M01_AXI_WSTRB          (io_PSmemory_2_1_wstrb),      
    .M01_AXI_WLAST          (io_PSmemory_2_1_wlast),      
    .M01_AXI_WVALID         (io_PSmemory_2_1_wvalid),    
    .M01_AXI_WREADY         (io_PSmemory_2_1_wready),   
    .M01_AXI_BID            (io_PSmemory_2_1_bid),         
    .M01_AXI_BRESP          (io_PSmemory_2_1_bresp),     
    .M01_AXI_BVALID         (io_PSmemory_2_1_bvalid),   
    .M01_AXI_BREADY         (io_PSmemory_2_1_bready),    
    .M01_AXI_ARID           (io_PSmemory_2_1_arid),        
    .M01_AXI_ARADDR         (io_PSmemory_2_1_araddr),    
    .M01_AXI_ARLEN          (io_PSmemory_2_1_arlen),      
    .M01_AXI_ARSIZE         (io_PSmemory_2_1_arsize),    
    .M01_AXI_ARBURST        (io_PSmemory_2_1_arburst),  
    .M01_AXI_ARLOCK         (io_PSmemory_2_1_arlock),    
    .M01_AXI_ARCACHE        (),                       
    .M01_AXI_ARPROT         (),                        
    .M01_AXI_ARVALID        (io_PSmemory_2_1_arvalid),  
    .M01_AXI_ARREADY        (io_PSmemory_2_1_arready), 
    .M01_AXI_RID            (io_PSmemory_2_1_rid),         
    .M01_AXI_RDATA          (io_PSmemory_2_1_rdata),     
    .M01_AXI_RRESP          (io_PSmemory_2_1_rresp),     
    .M01_AXI_RLAST          (io_PSmemory_2_1_rlast),     
    .M01_AXI_RVALID         (io_PSmemory_2_1_rvalid),   
    .M01_AXI_RREADY         (io_PSmemory_2_1_rready) 
    );
    
    wire [63:0]  io_PSmemory_3_0_awaddr;
    wire [5:0]   io_PSmemory_3_0_awid;
    wire [7:0]   io_PSmemory_3_0_awlen;
    wire [2:0]   io_PSmemory_3_0_awsize;
    wire [1:0]   io_PSmemory_3_0_awburst;
    wire         io_PSmemory_3_0_awlock;
    wire         io_PSmemory_3_0_awvalid;
    wire         io_PSmemory_3_0_awready;
    wire [63:0]  io_PSmemory_3_0_araddr;
    wire [5:0]   io_PSmemory_3_0_arid;
    wire [7:0]   io_PSmemory_3_0_arlen;
    wire [2:0]   io_PSmemory_3_0_arsize;
    wire [1:0]   io_PSmemory_3_0_arburst;
    wire         io_PSmemory_3_0_arlock;
    wire         io_PSmemory_3_0_arvalid;
    wire         io_PSmemory_3_0_arready;
    wire [511:0] io_PSmemory_3_0_wdata;
    wire [63:0]  io_PSmemory_3_0_wstrb;
    wire         io_PSmemory_3_0_wlast;
    wire         io_PSmemory_3_0_wvalid;
    wire         io_PSmemory_3_0_wready;
    wire  [511:0]io_PSmemory_3_0_rdata;
    wire  [5:0]  io_PSmemory_3_0_rid;
    wire         io_PSmemory_3_0_rlast;
    wire  [1:0]  io_PSmemory_3_0_rresp;
    wire         io_PSmemory_3_0_rvalid;
    wire         io_PSmemory_3_0_rready;
    wire  [1:0]  io_PSmemory_3_0_bresp;
    wire  [5:0]  io_PSmemory_3_0_bid;
    wire         io_PSmemory_3_0_bvalid;
    wire         io_PSmemory_3_0_bready;

    wire [63:0]  io_PSmemory_3_1_awaddr;
    wire [5:0]   io_PSmemory_3_1_awid;
    wire [7:0]   io_PSmemory_3_1_awlen;
    wire [2:0]   io_PSmemory_3_1_awsize;
    wire [1:0]   io_PSmemory_3_1_awburst;
    wire         io_PSmemory_3_1_awlock;
    wire         io_PSmemory_3_1_awvalid;
    wire         io_PSmemory_3_1_awready;
    wire [63:0]  io_PSmemory_3_1_araddr;
    wire [5:0]   io_PSmemory_3_1_arid;
    wire [7:0]   io_PSmemory_3_1_arlen;
    wire [2:0]   io_PSmemory_3_1_arsize;
    wire [1:0]   io_PSmemory_3_1_arburst;
    wire         io_PSmemory_3_1_arlock;
    wire         io_PSmemory_3_1_arvalid;
    wire         io_PSmemory_3_1_arready;
    wire [511:0] io_PSmemory_3_1_wdata;
    wire [63:0]  io_PSmemory_3_1_wstrb;
    wire         io_PSmemory_3_1_wlast;
    wire         io_PSmemory_3_1_wvalid;
    wire         io_PSmemory_3_1_wready;
    wire  [511:0]io_PSmemory_3_1_rdata;
    wire  [5:0]  io_PSmemory_3_1_rid;
    wire         io_PSmemory_3_1_rlast;
    wire  [1:0]  io_PSmemory_3_1_rresp;
    wire         io_PSmemory_3_1_rvalid;
    wire         io_PSmemory_3_1_rready;
    wire  [1:0]  io_PSmemory_3_1_bresp;
    wire  [5:0]  io_PSmemory_3_1_bid;
    wire         io_PSmemory_3_1_bvalid;
    wire         io_PSmemory_3_1_bready;

    memory u_hp3_memory(
    .gt_txusrclk(gt_txusrclk),
    .peripheral_reset(peripheral_reset),
    .M00_AXI_AWID           (io_PSmemory_3_0_awid),     
    .M00_AXI_AWADDR         (io_PSmemory_3_0_awaddr),   
    .M00_AXI_AWLEN          (io_PSmemory_3_0_awlen),    
    .M00_AXI_AWSIZE         (io_PSmemory_3_0_awsize),   
    .M00_AXI_AWBURST        (io_PSmemory_3_0_awburst),  
    .M00_AXI_AWLOCK         (io_PSmemory_3_0_awlock),   
    .M00_AXI_AWCACHE        (),  
    .M00_AXI_AWPROT         (),   
    .M00_AXI_AWVALID        (io_PSmemory_3_0_awvalid),  
    .M00_AXI_AWREADY        (io_PSmemory_3_0_awready), 
    .M00_AXI_WDATA          (io_PSmemory_3_0_wdata),    
    .M00_AXI_WSTRB          (io_PSmemory_3_0_wstrb),    
    .M00_AXI_WLAST          (io_PSmemory_3_0_wlast),    
    .M00_AXI_WVALID         (io_PSmemory_3_0_wvalid),   
    .M00_AXI_WREADY         (io_PSmemory_3_0_wready),  
    .M00_AXI_BID            (io_PSmemory_3_0_bid),     
    .M00_AXI_BRESP          (io_PSmemory_3_0_bresp),   
    .M00_AXI_BVALID         (io_PSmemory_3_0_bvalid),  
    .M00_AXI_BREADY         (io_PSmemory_3_0_bready),   
    .M00_AXI_ARID           (io_PSmemory_3_0_arid),     
    .M00_AXI_ARADDR         (io_PSmemory_3_0_araddr),   
    .M00_AXI_ARLEN          (io_PSmemory_3_0_arlen),    
    .M00_AXI_ARSIZE         (io_PSmemory_3_0_arsize),   
    .M00_AXI_ARBURST        (io_PSmemory_3_0_arburst),  
    .M00_AXI_ARLOCK         (io_PSmemory_3_0_arlock),   
    .M00_AXI_ARCACHE        (),  
    .M00_AXI_ARPROT         (),   
    .M00_AXI_ARVALID        (io_PSmemory_3_0_arvalid),  
    .M00_AXI_ARREADY        (io_PSmemory_3_0_arready), 
    .M00_AXI_RID            (io_PSmemory_3_0_rid),     
    .M00_AXI_RDATA          (io_PSmemory_3_0_rdata),   
    .M00_AXI_RRESP          (io_PSmemory_3_0_rresp),   
    .M00_AXI_RLAST          (io_PSmemory_3_0_rlast),   
    .M00_AXI_RVALID         (io_PSmemory_3_0_rvalid),  
    .M00_AXI_RREADY         (io_PSmemory_3_0_rready),   
                  
    .M01_AXI_AWID           (io_PSmemory_3_1_awid),        
    .M01_AXI_AWADDR         (io_PSmemory_3_1_awaddr),    
    .M01_AXI_AWLEN          (io_PSmemory_3_1_awlen),      
    .M01_AXI_AWSIZE         (io_PSmemory_3_1_awsize),    
    .M01_AXI_AWBURST        (io_PSmemory_3_1_awburst),  
    .M01_AXI_AWLOCK         (io_PSmemory_3_1_awlock),    
    .M01_AXI_AWCACHE        (),                       
    .M01_AXI_AWPROT         (),                        
    .M01_AXI_AWVALID        (io_PSmemory_3_1_awvalid),  
    .M01_AXI_AWREADY        (io_PSmemory_3_1_awready), 
    .M01_AXI_WDATA          (io_PSmemory_3_1_wdata),      
    .M01_AXI_WSTRB          (io_PSmemory_3_1_wstrb),      
    .M01_AXI_WLAST          (io_PSmemory_3_1_wlast),      
    .M01_AXI_WVALID         (io_PSmemory_3_1_wvalid),    
    .M01_AXI_WREADY         (io_PSmemory_3_1_wready),   
    .M01_AXI_BID            (io_PSmemory_3_1_bid),         
    .M01_AXI_BRESP          (io_PSmemory_3_1_bresp),     
    .M01_AXI_BVALID         (io_PSmemory_3_1_bvalid),   
    .M01_AXI_BREADY         (io_PSmemory_3_1_bready),    
    .M01_AXI_ARID           (io_PSmemory_3_1_arid),        
    .M01_AXI_ARADDR         (io_PSmemory_3_1_araddr),    
    .M01_AXI_ARLEN          (io_PSmemory_3_1_arlen),      
    .M01_AXI_ARSIZE         (io_PSmemory_3_1_arsize),    
    .M01_AXI_ARBURST        (io_PSmemory_3_1_arburst),  
    .M01_AXI_ARLOCK         (io_PSmemory_3_1_arlock),    
    .M01_AXI_ARCACHE        (),                       
    .M01_AXI_ARPROT         (),                        
    .M01_AXI_ARVALID        (io_PSmemory_3_1_arvalid),  
    .M01_AXI_ARREADY        (io_PSmemory_3_1_arready), 
    .M01_AXI_RID            (io_PSmemory_3_1_rid),         
    .M01_AXI_RDATA          (io_PSmemory_3_1_rdata),     
    .M01_AXI_RRESP          (io_PSmemory_3_1_rresp),     
    .M01_AXI_RLAST          (io_PSmemory_3_1_rlast),     
    .M01_AXI_RVALID         (io_PSmemory_3_1_rvalid),   
    .M01_AXI_RREADY         (io_PSmemory_3_1_rready) 
    );
     
  wire [63:0]  io_PLmemory_0_awaddr;
    wire [5:0]   io_PLmemory_0_awid;
    wire [7:0]   io_PLmemory_0_awlen;
    wire [2:0]   io_PLmemory_0_awsize;
    wire [1:0]   io_PLmemory_0_awburst;
    wire         io_PLmemory_0_awlock;
    wire         io_PLmemory_0_awvalid;
    wire         io_PLmemory_0_awready;
    wire [63:0]  io_PLmemory_0_araddr;
    wire [5:0]   io_PLmemory_0_arid;
    wire [7:0]   io_PLmemory_0_arlen;
    wire [2:0]   io_PLmemory_0_arsize;
    wire [1:0]   io_PLmemory_0_arburst;
    wire         io_PLmemory_0_arlock;
    wire         io_PLmemory_0_arvalid;
    wire         io_PLmemory_0_arready;
    wire [511:0] io_PLmemory_0_wdata;
    wire [63:0]  io_PLmemory_0_wstrb;
    wire         io_PLmemory_0_wlast;
    wire         io_PLmemory_0_wvalid;
    wire         io_PLmemory_0_wready;
    wire  [511:0]io_PLmemory_0_rdata;
    wire  [5:0]  io_PLmemory_0_rid;
    wire         io_PLmemory_0_rlast;
    wire  [1:0]  io_PLmemory_0_rresp;
    wire         io_PLmemory_0_rvalid;
    wire         io_PLmemory_0_rready;
    wire  [1:0]  io_PLmemory_0_bresp;
    wire  [5:0]  io_PLmemory_0_bid;
    wire         io_PLmemory_0_bvalid;
    wire         io_PLmemory_0_bready;

    wire [63:0]  io_PLmemory_1_awaddr;
    wire [5:0]   io_PLmemory_1_awid;
    wire [7:0]   io_PLmemory_1_awlen;
    wire [2:0]   io_PLmemory_1_awsize;
    wire [1:0]   io_PLmemory_1_awburst;
    wire         io_PLmemory_1_awlock;
    wire         io_PLmemory_1_awvalid;
    wire         io_PLmemory_1_awready;
    wire [63:0]  io_PLmemory_1_araddr;
    wire [5:0]   io_PLmemory_1_arid;
    wire [7:0]   io_PLmemory_1_arlen;
    wire [2:0]   io_PLmemory_1_arsize;
    wire [1:0]   io_PLmemory_1_arburst;
    wire         io_PLmemory_1_arlock;
    wire         io_PLmemory_1_arvalid;
    wire         io_PLmemory_1_arready;
    wire [511:0] io_PLmemory_1_wdata;
    wire [63:0]  io_PLmemory_1_wstrb;
    wire         io_PLmemory_1_wlast;
    wire         io_PLmemory_1_wvalid;
    wire         io_PLmemory_1_wready;
    wire  [511:0]io_PLmemory_1_rdata;
    wire  [5:0]  io_PLmemory_1_rid;
    wire         io_PLmemory_1_rlast;
    wire  [1:0]  io_PLmemory_1_rresp;
    wire         io_PLmemory_1_rvalid;
    wire         io_PLmemory_1_rready;
    wire  [1:0]  io_PLmemory_1_bresp;
    wire  [5:0]  io_PLmemory_1_bid;
    wire         io_PLmemory_1_bvalid;
    wire         io_PLmemory_1_bready;
  
  wire         io_PSmempory_aw_ready;
  wire         io_PSmempory_aw_valid;
  wire [63:0]  io_PSmempory_aw_bits_awaddr;
  wire [5:0]   io_PSmempory_aw_bits_awid;
  wire [7:0]   io_PSmempory_aw_bits_awlen;
  wire [2:0]   io_PSmempory_aw_bits_awsize;
  wire [1:0]   io_PSmempory_aw_bits_awburst;
  wire         io_PSmempory_aw_bits_awlock;
  wire         io_PSmempory_ar_ready;
  wire         io_PSmempory_ar_valid;
  wire [63:0]  io_PSmempory_ar_bits_araddr;
  wire [5:0]   io_PSmempory_ar_bits_arid;
  wire [7:0]   io_PSmempory_ar_bits_arlen;
  wire [2:0]   io_PSmempory_ar_bits_arsize;
  wire [1:0]   io_PSmempory_ar_bits_arburst;
  wire         io_PSmempory_ar_bits_arlock;
  wire         io_PSmempory_w_ready;
  wire         io_PSmempory_w_valid;
  wire [127:0] io_PSmempory_w_bits_wdata;
  wire [15:0]  io_PSmempory_w_bits_wstrb;
  wire         io_PSmempory_w_bits_wlast;
  wire         io_PSmempory_r_ready;
  wire         io_PSmempory_r_valid;
  wire [127:0] io_PSmempory_r_bits_rdata;
  wire [5:0]   io_PSmempory_r_bits_rid;
  wire         io_PSmempory_r_bits_rlast;
  wire         io_PSmempory_b_ready;
  wire         io_PSmempory_b_valid;
  wire [1:0]   io_PSmempory_b_bits_bresp;
  wire [5:0]   io_PSmempory_b_bits_bid;

  wire         io_PSmempory_1_aw_ready;
  wire         io_PSmempory_1_aw_valid;
  wire [63:0]  io_PSmempory_1_aw_bits_awaddr;
  wire [5:0]   io_PSmempory_1_aw_bits_awid;
  wire [7:0]   io_PSmempory_1_aw_bits_awlen;
  wire [2:0]   io_PSmempory_1_aw_bits_awsize;
  wire [1:0]   io_PSmempory_1_aw_bits_awburst;
  wire         io_PSmempory_1_aw_bits_awlock;
  wire         io_PSmempory_1_ar_ready;
  wire         io_PSmempory_1_ar_valid;
  wire [63:0]  io_PSmempory_1_ar_bits_araddr;
  wire [5:0]   io_PSmempory_1_ar_bits_arid;
  wire [7:0]   io_PSmempory_1_ar_bits_arlen;
  wire [2:0]   io_PSmempory_1_ar_bits_arsize;
  wire [1:0]   io_PSmempory_1_ar_bits_arburst;
  wire         io_PSmempory_1_ar_bits_arlock;
  wire         io_PSmempory_1_w_ready;
  wire         io_PSmempory_1_w_valid;
  wire [127:0] io_PSmempory_1_w_bits_wdata;
  wire [15:0]  io_PSmempory_1_w_bits_wstrb;
  wire         io_PSmempory_1_w_bits_wlast;
  wire         io_PSmempory_1_r_ready;
  wire         io_PSmempory_1_r_valid;
  wire [127:0] io_PSmempory_1_r_bits_rdata;
  wire [5:0]   io_PSmempory_1_r_bits_rid;
  wire         io_PSmempory_1_r_bits_rlast;
  wire         io_PSmempory_1_b_ready;
  wire         io_PSmempory_1_b_valid;
  wire [1:0]   io_PSmempory_1_b_bits_bresp;
  wire [5:0]   io_PSmempory_1_b_bits_bid;

  wire         io_PSmempory_2_aw_ready;
  wire         io_PSmempory_2_aw_valid;
  wire [63:0]  io_PSmempory_2_aw_bits_awaddr;
  wire [5:0]   io_PSmempory_2_aw_bits_awid;
  wire [7:0]   io_PSmempory_2_aw_bits_awlen;
  wire [2:0]   io_PSmempory_2_aw_bits_awsize;
  wire [1:0]   io_PSmempory_2_aw_bits_awburst;
  wire         io_PSmempory_2_aw_bits_awlock;
  wire         io_PSmempory_2_ar_ready;
  wire         io_PSmempory_2_ar_valid;
  wire [63:0]  io_PSmempory_2_ar_bits_araddr;
  wire [5:0]   io_PSmempory_2_ar_bits_arid;
  wire [7:0]   io_PSmempory_2_ar_bits_arlen;
  wire [2:0]   io_PSmempory_2_ar_bits_arsize;
  wire [1:0]   io_PSmempory_2_ar_bits_arburst;
  wire         io_PSmempory_2_ar_bits_arlock;
  wire         io_PSmempory_2_w_ready;
  wire         io_PSmempory_2_w_valid;
  wire [127:0] io_PSmempory_2_w_bits_wdata;
  wire [15:0]  io_PSmempory_2_w_bits_wstrb;
  wire         io_PSmempory_2_w_bits_wlast;
  wire         io_PSmempory_2_r_ready;
  wire         io_PSmempory_2_r_valid;
  wire [127:0] io_PSmempory_2_r_bits_rdata;
  wire [5:0]   io_PSmempory_2_r_bits_rid;
  wire         io_PSmempory_2_r_bits_rlast;
  wire         io_PSmempory_2_b_ready;
  wire         io_PSmempory_2_b_valid;
  wire [1:0]   io_PSmempory_2_b_bits_bresp;
  wire [5:0]   io_PSmempory_2_b_bits_bid;

  wire         io_PSmempory_3_aw_ready;
  wire         io_PSmempory_3_aw_valid;
  wire [63:0]  io_PSmempory_3_aw_bits_awaddr;
  wire [5:0]   io_PSmempory_3_aw_bits_awid;
  wire [7:0]   io_PSmempory_3_aw_bits_awlen;
  wire [2:0]   io_PSmempory_3_aw_bits_awsize;
  wire [1:0]   io_PSmempory_3_aw_bits_awburst;
  wire         io_PSmempory_3_aw_bits_awlock;
  wire         io_PSmempory_3_ar_ready;
  wire         io_PSmempory_3_ar_valid;
  wire [63:0]  io_PSmempory_3_ar_bits_araddr;
  wire [5:0]   io_PSmempory_3_ar_bits_arid;
  wire [7:0]   io_PSmempory_3_ar_bits_arlen;
  wire [2:0]   io_PSmempory_3_ar_bits_arsize;
  wire [1:0]   io_PSmempory_3_ar_bits_arburst;
  wire         io_PSmempory_3_ar_bits_arlock;
  wire         io_PSmempory_3_w_ready;
  wire         io_PSmempory_3_w_valid;
  wire [127:0] io_PSmempory_3_w_bits_wdata;
  wire [15:0]  io_PSmempory_3_w_bits_wstrb;
  wire         io_PSmempory_3_w_bits_wlast;
  wire         io_PSmempory_3_r_ready;
  wire         io_PSmempory_3_r_valid;
  wire [127:0] io_PSmempory_3_r_bits_rdata;
  wire [5:0]   io_PSmempory_3_r_bits_rid;
  wire         io_PSmempory_3_r_bits_rlast;
  wire         io_PSmempory_3_b_ready;
  wire         io_PSmempory_3_b_valid;
  wire [1:0]   io_PSmempory_3_b_bits_bresp;
  wire [5:0]   io_PSmempory_3_b_bits_bid;

  wire         io_Re_memory_out_aw_ready;
  wire         io_Re_memory_out_aw_valid;
  wire [63:0]  io_Re_memory_out_aw_bits_awaddr;
  wire [5:0]   io_Re_memory_out_aw_bits_awid;
  wire [7:0]   io_Re_memory_out_aw_bits_awlen;
  wire [2:0]   io_Re_memory_out_aw_bits_awsize;
  wire [1:0]   io_Re_memory_out_aw_bits_awburst;
  wire         io_Re_memory_out_aw_bits_awlock;
  wire         io_Re_memory_out_ar_ready;
  wire         io_Re_memory_out_ar_valid;
  wire [63:0]  io_Re_memory_out_ar_bits_araddr;
  wire [5:0]   io_Re_memory_out_ar_bits_arid;
  wire [7:0]   io_Re_memory_out_ar_bits_arlen;
  wire [2:0]   io_Re_memory_out_ar_bits_arsize;
  wire [1:0]   io_Re_memory_out_ar_bits_arburst;
  wire         io_Re_memory_out_ar_bits_arlock;
  wire         io_Re_memory_out_w_ready;
  wire         io_Re_memory_out_w_valid;
  wire [511:0] io_Re_memory_out_w_bits_wdata;
  wire [63:0]  io_Re_memory_out_w_bits_wstrb;
  wire         io_Re_memory_out_w_bits_wlast;
  wire         io_Re_memory_out_r_ready;
  wire         io_Re_memory_out_r_valid;
  wire [511:0] io_Re_memory_out_r_bits_rdata;
  wire [5:0]   io_Re_memory_out_r_bits_rid;
  wire         io_Re_memory_out_r_bits_rlast;
  wire         io_Re_memory_out_b_ready;
  wire         io_Re_memory_out_b_valid;
  wire [1:0]   io_Re_memory_out_b_bits_bresp;
  wire [5:0]   io_Re_memory_out_b_bits_bid;

  wire         io_Re_memory_in_aw_ready;
  wire         io_Re_memory_in_aw_valid;
  wire [63:0]  io_Re_memory_in_aw_bits_awaddr;
  wire [9:0]   io_Re_memory_in_aw_bits_awid;
  wire [7:0]   io_Re_memory_in_aw_bits_awlen;
  wire [2:0]   io_Re_memory_in_aw_bits_awsize;
  wire [1:0]   io_Re_memory_in_aw_bits_awburst;
  wire         io_Re_memory_in_aw_bits_awlock;
  wire         io_Re_memory_in_ar_ready;
  wire         io_Re_memory_in_ar_valid;
  wire [63:0]  io_Re_memory_in_ar_bits_araddr;
  wire [9:0]   io_Re_memory_in_ar_bits_arid;
  wire [7:0]   io_Re_memory_in_ar_bits_arlen;
  wire [2:0]   io_Re_memory_in_ar_bits_arsize;
  wire [1:0]   io_Re_memory_in_ar_bits_arburst;
  wire         io_Re_memory_in_ar_bits_arlock;
  wire         io_Re_memory_in_w_ready;
  wire         io_Re_memory_in_w_valid;
  wire [511:0] io_Re_memory_in_w_bits_wdata;
  wire [63:0]  io_Re_memory_in_w_bits_wstrb;
  wire         io_Re_memory_in_w_bits_wlast;
  wire         io_Re_memory_in_r_ready;
  wire         io_Re_memory_in_r_valid;
  wire [511:0] io_Re_memory_in_r_bits_rdata;
  wire [9:0]   io_Re_memory_in_r_bits_rid;
  wire         io_Re_memory_in_r_bits_rlast;
  wire         io_Re_memory_in_b_ready;
  wire         io_Re_memory_in_b_valid;
  wire [1:0]   io_Re_memory_in_b_bits_bresp;
  wire [9:0]   io_Re_memory_in_b_bits_bid;

  wire [63:0]  bfs_io_config_awaddr;
  wire         bfs_io_config_awvalid;
  wire         bfs_io_config_awready;
  wire [63:0]  bfs_io_config_araddr;
  wire         bfs_io_config_arvalid;
  wire         bfs_io_config_arready;
  wire [31:0]  bfs_io_config_wdata;
  wire [3:0]   bfs_io_config_wstrb;
  wire         bfs_io_config_wvalid;
  wire         bfs_io_config_wready;
  wire [31:0]  bfs_io_config_rdata;
  wire [1:0]   bfs_io_config_rresp;
  wire         bfs_io_config_rvalid;
  wire         bfs_io_config_rready;
  wire [1:0]   bfs_io_config_bresp;
  wire         bfs_io_config_bvalid;
  wire         bfs_io_config_bready;

    design_1 u_xbar(
      .INTERCONNECT_ACLK      (gt_txusrclk),
      .INTERCONNECT_ARESETN   (~peripheral_reset),
      .clk_doce                 (doceclk),
      .doce_resetn              (~peripheral_reset),
      .clk_cmac                  (cmacclk),
      .cmac_resetn              (~peripheral_reset),

      .doce_axis_rxd_tdata    (doce_axis_rxd_tdata),
      .doce_axis_rxd_tkeep    (doce_axis_rxd_tkeep),
      .doce_axis_rxd_tlast    (doce_axis_rxd_tlast),
      .doce_axis_rxd_tready   (doce_axis_rxd_tready),
      .doce_axis_rxd_tvalid   (doce_axis_rxd_tvalid),
      .doce_axis_txd_tdata    (doce_axis_txd_tdata),
      .doce_axis_txd_tkeep    (doce_axis_txd_tkeep),
      .doce_axis_txd_tlast    (doce_axis_txd_tlast),
      .doce_axis_txd_tready   (doce_axis_txd_tready),
      .doce_axis_txd_tvalid   (doce_axis_txd_tvalid),

      .io_PLmemory_0_awid           ({1'b0, io_PLmemory_0_awid[5:0]}),
      .io_PLmemory_0_awaddr         (io_PLmemory_0_awaddr),
      .io_PLmemory_0_awlen          (io_PLmemory_0_awlen),
      .io_PLmemory_0_awsize         (io_PLmemory_0_awsize),
      .io_PLmemory_0_awburst        (io_PLmemory_0_awburst),
      .io_PLmemory_0_awlock         (io_PLmemory_0_awlock),
      .io_PLmemory_0_awvalid        (io_PLmemory_0_awvalid),
      .io_PLmemory_0_awready        (io_PLmemory_0_awready),
      .io_PLmemory_0_wdata          (io_PLmemory_0_wdata),
      .io_PLmemory_0_wstrb          (io_PLmemory_0_wstrb),
      .io_PLmemory_0_wlast          (io_PLmemory_0_wlast),
      .io_PLmemory_0_wvalid         (io_PLmemory_0_wvalid),
      .io_PLmemory_0_wready         (io_PLmemory_0_wready),
      .io_PLmemory_0_bid            (io_PLmemory_0_bid),
      .io_PLmemory_0_bresp          (io_PLmemory_0_bresp),
      .io_PLmemory_0_bvalid         (io_PLmemory_0_bvalid),
      .io_PLmemory_0_bready         (io_PLmemory_0_bready),
      .io_PLmemory_0_arid           ({1'b0, io_PLmemory_0_arid[5:0]}),
      .io_PLmemory_0_araddr         (io_PLmemory_0_araddr),
      .io_PLmemory_0_arlen          (io_PLmemory_0_arlen),
      .io_PLmemory_0_arsize         (io_PLmemory_0_arsize),
      .io_PLmemory_0_arburst        (io_PLmemory_0_arburst),
      .io_PLmemory_0_arlock         (io_PLmemory_0_arlock),
      .io_PLmemory_0_arvalid        (io_PLmemory_0_arvalid),
      .io_PLmemory_0_arready        (io_PLmemory_0_arready),
      .io_PLmemory_0_rid            (io_PLmemory_0_rid),
      .io_PLmemory_0_rdata          (io_PLmemory_0_rdata),
      .io_PLmemory_0_rresp          (io_PLmemory_0_rresp),
      .io_PLmemory_0_rlast          (io_PLmemory_0_rlast),
      .io_PLmemory_0_rvalid         (io_PLmemory_0_rvalid),
      .io_PLmemory_0_rready         (io_PLmemory_0_rready),

      .io_PLmemory_1_awid           ({1'b0, io_PLmemory_1_awid[5:0]}),
      .io_PLmemory_1_awaddr         (io_PLmemory_1_awaddr),
      .io_PLmemory_1_awlen          (io_PLmemory_1_awlen),
      .io_PLmemory_1_awsize         (io_PLmemory_1_awsize),
      .io_PLmemory_1_awburst        (io_PLmemory_1_awburst),
      .io_PLmemory_1_awlock         (io_PLmemory_1_awlock),
      .io_PLmemory_1_awvalid        (io_PLmemory_1_awvalid),
      .io_PLmemory_1_awready        (io_PLmemory_1_awready),
      .io_PLmemory_1_wdata          (io_PLmemory_1_wdata),
      .io_PLmemory_1_wstrb          (io_PLmemory_1_wstrb),
      .io_PLmemory_1_wlast          (io_PLmemory_1_wlast),
      .io_PLmemory_1_wvalid         (io_PLmemory_1_wvalid),
      .io_PLmemory_1_wready         (io_PLmemory_1_wready),
      .io_PLmemory_1_bid            (io_PLmemory_1_bid),
      .io_PLmemory_1_bresp          (io_PLmemory_1_bresp),
      .io_PLmemory_1_bvalid         (io_PLmemory_1_bvalid),
      .io_PLmemory_1_bready         (io_PLmemory_1_bready),
      .io_PLmemory_1_arid           ({1'b0, io_PLmemory_1_arid[5:0]}),
      .io_PLmemory_1_araddr         (io_PLmemory_1_araddr),
      .io_PLmemory_1_arlen          (io_PLmemory_1_arlen),
      .io_PLmemory_1_arsize         (io_PLmemory_1_arsize),
      .io_PLmemory_1_arburst        (io_PLmemory_1_arburst),
      .io_PLmemory_1_arlock         (io_PLmemory_1_arlock),
      .io_PLmemory_1_arvalid        (io_PLmemory_1_arvalid),
      .io_PLmemory_1_arready        (io_PLmemory_1_arready),
      .io_PLmemory_1_rid            (io_PLmemory_1_rid),
      .io_PLmemory_1_rdata          (io_PLmemory_1_rdata),
      .io_PLmemory_1_rresp          (io_PLmemory_1_rresp),
      .io_PLmemory_1_rlast          (io_PLmemory_1_rlast),
      .io_PLmemory_1_rvalid         (io_PLmemory_1_rvalid),
      .io_PLmemory_1_rready         (io_PLmemory_1_rready),

      //.io_PLmemory_awid           (io_PLmemory_awid),
      .io_PLmemory_awaddr         (io_PLmemory_awaddr),
      .io_PLmemory_awlen          (io_PLmemory_awlen),
      .io_PLmemory_awsize         (io_PLmemory_awsize),
      .io_PLmemory_awburst        (io_PLmemory_awburst),
      .io_PLmemory_awlock         (io_PLmemory_awlock),
      .io_PLmemory_awvalid        (io_PLmemory_awvalid),
      .io_PLmemory_awready        (io_PLmemory_awready),
      .io_PLmemory_wdata          (io_PLmemory_wdata),
      .io_PLmemory_wstrb          (io_PLmemory_wstrb),
      .io_PLmemory_wlast          (io_PLmemory_wlast),
      .io_PLmemory_wvalid         (io_PLmemory_wvalid),
      .io_PLmemory_wready         (io_PLmemory_wready),
      //.io_PLmemory_bid            (io_PLmemory_bid),
      .io_PLmemory_bresp          (io_PLmemory_bresp),
      .io_PLmemory_bvalid         (io_PLmemory_bvalid),
      .io_PLmemory_bready         (io_PLmemory_bready),
      //.io_PLmemory_arid           (io_PLmemory_arid),
      .io_PLmemory_araddr         (io_PLmemory_araddr),
      .io_PLmemory_arlen          (io_PLmemory_arlen),
      .io_PLmemory_arsize         (io_PLmemory_arsize),
      .io_PLmemory_arburst        (io_PLmemory_arburst),
      .io_PLmemory_arlock         (io_PLmemory_arlock),
      .io_PLmemory_arvalid        (io_PLmemory_arvalid),
      .io_PLmemory_arready        (io_PLmemory_arready),
      //.io_PLmemory_rid            (io_PLmemory_rid),
      .io_PLmemory_rdata          (io_PLmemory_rdata),
      .io_PLmemory_rresp          (io_PLmemory_rresp),
      .io_PLmemory_rlast          (io_PLmemory_rlast),
      .io_PLmemory_rvalid         (io_PLmemory_rvalid),
      .io_PLmemory_rready         (io_PLmemory_rready),
      
      //.io_PSmemory_0_0_awid           (io_PSmemory_0_0_awid),
      .io_PSmemory_0_0_awaddr         (io_PSmemory_0_0_awaddr),
      .io_PSmemory_0_0_awlen          (io_PSmemory_0_0_awlen),
      .io_PSmemory_0_0_awsize         (io_PSmemory_0_0_awsize),
      .io_PSmemory_0_0_awburst        (io_PSmemory_0_0_awburst),
      .io_PSmemory_0_0_awlock         (io_PSmemory_0_0_awlock),
      .io_PSmemory_0_0_awvalid        (io_PSmemory_0_0_awvalid),
      .io_PSmemory_0_0_awready        (io_PSmemory_0_0_awready),
      .io_PSmemory_0_0_wdata          (io_PSmemory_0_0_wdata),
      .io_PSmemory_0_0_wstrb          (io_PSmemory_0_0_wstrb),
      .io_PSmemory_0_0_wlast          (io_PSmemory_0_0_wlast),
      .io_PSmemory_0_0_wvalid         (io_PSmemory_0_0_wvalid),
      .io_PSmemory_0_0_wready         (io_PSmemory_0_0_wready),
      //.io_PSmemory_0_0_bid            (io_PSmemory_0_0_bid),
      .io_PSmemory_0_0_bresp          (io_PSmemory_0_0_bresp),
      .io_PSmemory_0_0_bvalid         (io_PSmemory_0_0_bvalid),
      .io_PSmemory_0_0_bready         (io_PSmemory_0_0_bready),
      //.io_PSmemory_0_0_arid           (io_PSmemory_0_0_arid),
      .io_PSmemory_0_0_araddr         (io_PSmemory_0_0_araddr),
      .io_PSmemory_0_0_arlen          (io_PSmemory_0_0_arlen),
      .io_PSmemory_0_0_arsize         (io_PSmemory_0_0_arsize),
      .io_PSmemory_0_0_arburst        (io_PSmemory_0_0_arburst),
      .io_PSmemory_0_0_arlock         (io_PSmemory_0_0_arlock),
      .io_PSmemory_0_0_arvalid        (io_PSmemory_0_0_arvalid),
      .io_PSmemory_0_0_arready        (io_PSmemory_0_0_arready),
      //.io_PSmemory_0_0_rid            (io_PSmemory_0_0_rid),
      .io_PSmemory_0_0_rdata          (io_PSmemory_0_0_rdata),
      .io_PSmemory_0_0_rresp          (io_PSmemory_0_0_rresp),
      .io_PSmemory_0_0_rlast          (io_PSmemory_0_0_rlast),
      .io_PSmemory_0_0_rvalid         (io_PSmemory_0_0_rvalid),
      .io_PSmemory_0_0_rready         (io_PSmemory_0_0_rready),
      
      //.io_PSmemory_0_1_awid           (io_PSmemory_0_1_awid),
      .io_PSmemory_0_1_awaddr         (io_PSmemory_0_1_awaddr),
      .io_PSmemory_0_1_awlen          (io_PSmemory_0_1_awlen),
      .io_PSmemory_0_1_awsize         (io_PSmemory_0_1_awsize),
      .io_PSmemory_0_1_awburst        (io_PSmemory_0_1_awburst),
      .io_PSmemory_0_1_awlock         (io_PSmemory_0_1_awlock),
      .io_PSmemory_0_1_awvalid        (io_PSmemory_0_1_awvalid),
      .io_PSmemory_0_1_awready        (io_PSmemory_0_1_awready),
      .io_PSmemory_0_1_wdata          (io_PSmemory_0_1_wdata),
      .io_PSmemory_0_1_wstrb          (io_PSmemory_0_1_wstrb),
      .io_PSmemory_0_1_wlast          (io_PSmemory_0_1_wlast),
      .io_PSmemory_0_1_wvalid         (io_PSmemory_0_1_wvalid),
      .io_PSmemory_0_1_wready         (io_PSmemory_0_1_wready),
      //.io_PSmemory_0_1_bid            (io_PSmemory_0_1_bid),
      .io_PSmemory_0_1_bresp          (io_PSmemory_0_1_bresp),
      .io_PSmemory_0_1_bvalid         (io_PSmemory_0_1_bvalid),
      .io_PSmemory_0_1_bready         (io_PSmemory_0_1_bready),
      //.io_PSmemory_0_1_arid           (io_PSmemory_0_1_arid),
      .io_PSmemory_0_1_araddr         (io_PSmemory_0_1_araddr),
      .io_PSmemory_0_1_arlen          (io_PSmemory_0_1_arlen),
      .io_PSmemory_0_1_arsize         (io_PSmemory_0_1_arsize),
      .io_PSmemory_0_1_arburst        (io_PSmemory_0_1_arburst),
      .io_PSmemory_0_1_arlock         (io_PSmemory_0_1_arlock),
      .io_PSmemory_0_1_arvalid        (io_PSmemory_0_1_arvalid),
      .io_PSmemory_0_1_arready        (io_PSmemory_0_1_arready),
      //.io_PSmemory_0_1_rid            (io_PSmemory_0_1_rid),
      .io_PSmemory_0_1_rdata          (io_PSmemory_0_1_rdata),
      .io_PSmemory_0_1_rresp          (io_PSmemory_0_1_rresp),
      .io_PSmemory_0_1_rlast          (io_PSmemory_0_1_rlast),
      .io_PSmemory_0_1_rvalid         (io_PSmemory_0_1_rvalid),
      .io_PSmemory_0_1_rready         (io_PSmemory_0_1_rready),
      
      //.io_PSmemory_1_0_awid           (io_PSmemory_1_0_awid),
      .io_PSmemory_1_0_awaddr         (io_PSmemory_1_0_awaddr),
      .io_PSmemory_1_0_awlen          (io_PSmemory_1_0_awlen),
      .io_PSmemory_1_0_awsize         (io_PSmemory_1_0_awsize),
      .io_PSmemory_1_0_awburst        (io_PSmemory_1_0_awburst),
      .io_PSmemory_1_0_awlock         (io_PSmemory_1_0_awlock),
      .io_PSmemory_1_0_awvalid        (io_PSmemory_1_0_awvalid),
      .io_PSmemory_1_0_awready        (io_PSmemory_1_0_awready),
      .io_PSmemory_1_0_wdata          (io_PSmemory_1_0_wdata),
      .io_PSmemory_1_0_wstrb          (io_PSmemory_1_0_wstrb),
      .io_PSmemory_1_0_wlast          (io_PSmemory_1_0_wlast),
      .io_PSmemory_1_0_wvalid         (io_PSmemory_1_0_wvalid),
      .io_PSmemory_1_0_wready         (io_PSmemory_1_0_wready),
      //.io_PSmemory_1_0_bid            (io_PSmemory_1_0_bid),
      .io_PSmemory_1_0_bresp          (io_PSmemory_1_0_bresp),
      .io_PSmemory_1_0_bvalid         (io_PSmemory_1_0_bvalid),
      .io_PSmemory_1_0_bready         (io_PSmemory_1_0_bready),
      //.io_PSmemory_1_0_arid           (io_PSmemory_1_0_arid),
      .io_PSmemory_1_0_araddr         (io_PSmemory_1_0_araddr),
      .io_PSmemory_1_0_arlen          (io_PSmemory_1_0_arlen),
      .io_PSmemory_1_0_arsize         (io_PSmemory_1_0_arsize),
      .io_PSmemory_1_0_arburst        (io_PSmemory_1_0_arburst),
      .io_PSmemory_1_0_arlock         (io_PSmemory_1_0_arlock),
      .io_PSmemory_1_0_arvalid        (io_PSmemory_1_0_arvalid),
      .io_PSmemory_1_0_arready        (io_PSmemory_1_0_arready),
      //.io_PSmemory_1_0_rid            (io_PSmemory_1_0_rid),
      .io_PSmemory_1_0_rdata          (io_PSmemory_1_0_rdata),
      .io_PSmemory_1_0_rresp          (io_PSmemory_1_0_rresp),
      .io_PSmemory_1_0_rlast          (io_PSmemory_1_0_rlast),
      .io_PSmemory_1_0_rvalid         (io_PSmemory_1_0_rvalid),
      .io_PSmemory_1_0_rready         (io_PSmemory_1_0_rready),
      
      //.io_PSmemory_1_1_awid           (io_PSmemory_1_1_awid),
      .io_PSmemory_1_1_awaddr         (io_PSmemory_1_1_awaddr),
      .io_PSmemory_1_1_awlen          (io_PSmemory_1_1_awlen),
      .io_PSmemory_1_1_awsize         (io_PSmemory_1_1_awsize),
      .io_PSmemory_1_1_awburst        (io_PSmemory_1_1_awburst),
      .io_PSmemory_1_1_awlock         (io_PSmemory_1_1_awlock),
      .io_PSmemory_1_1_awvalid        (io_PSmemory_1_1_awvalid),
      .io_PSmemory_1_1_awready        (io_PSmemory_1_1_awready),
      .io_PSmemory_1_1_wdata          (io_PSmemory_1_1_wdata),
      .io_PSmemory_1_1_wstrb          (io_PSmemory_1_1_wstrb),
      .io_PSmemory_1_1_wlast          (io_PSmemory_1_1_wlast),
      .io_PSmemory_1_1_wvalid         (io_PSmemory_1_1_wvalid),
      .io_PSmemory_1_1_wready         (io_PSmemory_1_1_wready),
      //.io_PSmemory_1_1_bid            (io_PSmemory_1_1_bid),
      .io_PSmemory_1_1_bresp          (io_PSmemory_1_1_bresp),
      .io_PSmemory_1_1_bvalid         (io_PSmemory_1_1_bvalid),
      .io_PSmemory_1_1_bready         (io_PSmemory_1_1_bready),
      //.io_PSmemory_1_1_arid           (io_PSmemory_1_1_arid),
      .io_PSmemory_1_1_araddr         (io_PSmemory_1_1_araddr),
      .io_PSmemory_1_1_arlen          (io_PSmemory_1_1_arlen),
      .io_PSmemory_1_1_arsize         (io_PSmemory_1_1_arsize),
      .io_PSmemory_1_1_arburst        (io_PSmemory_1_1_arburst),
      .io_PSmemory_1_1_arlock         (io_PSmemory_1_1_arlock),
      .io_PSmemory_1_1_arvalid        (io_PSmemory_1_1_arvalid),
      .io_PSmemory_1_1_arready        (io_PSmemory_1_1_arready),
      //.io_PSmemory_1_1_rid            (io_PSmemory_1_1_rid),
      .io_PSmemory_1_1_rdata          (io_PSmemory_1_1_rdata),
      .io_PSmemory_1_1_rresp          (io_PSmemory_1_1_rresp),
      .io_PSmemory_1_1_rlast          (io_PSmemory_1_1_rlast),
      .io_PSmemory_1_1_rvalid         (io_PSmemory_1_1_rvalid),
      .io_PSmemory_1_1_rready         (io_PSmemory_1_1_rready),
      
      //.io_PSmemory_2_0_awid           (io_PSmemory_2_0_awid),
      .io_PSmemory_2_0_awaddr         (io_PSmemory_2_0_awaddr),
      .io_PSmemory_2_0_awlen          (io_PSmemory_2_0_awlen),
      .io_PSmemory_2_0_awsize         (io_PSmemory_2_0_awsize),
      .io_PSmemory_2_0_awburst        (io_PSmemory_2_0_awburst),
      .io_PSmemory_2_0_awlock         (io_PSmemory_2_0_awlock),
      .io_PSmemory_2_0_awvalid        (io_PSmemory_2_0_awvalid),
      .io_PSmemory_2_0_awready        (io_PSmemory_2_0_awready),
      .io_PSmemory_2_0_wdata          (io_PSmemory_2_0_wdata),
      .io_PSmemory_2_0_wstrb          (io_PSmemory_2_0_wstrb),
      .io_PSmemory_2_0_wlast          (io_PSmemory_2_0_wlast),
      .io_PSmemory_2_0_wvalid         (io_PSmemory_2_0_wvalid),
      .io_PSmemory_2_0_wready         (io_PSmemory_2_0_wready),
      //.io_PSmemory_2_0_bid            (io_PSmemory_2_0_bid),
      .io_PSmemory_2_0_bresp          (io_PSmemory_2_0_bresp),
      .io_PSmemory_2_0_bvalid         (io_PSmemory_2_0_bvalid),
      .io_PSmemory_2_0_bready         (io_PSmemory_2_0_bready),
      //.io_PSmemory_2_0_arid           (io_PSmemory_2_0_arid),
      .io_PSmemory_2_0_araddr         (io_PSmemory_2_0_araddr),
      .io_PSmemory_2_0_arlen          (io_PSmemory_2_0_arlen),
      .io_PSmemory_2_0_arsize         (io_PSmemory_2_0_arsize),
      .io_PSmemory_2_0_arburst        (io_PSmemory_2_0_arburst),
      .io_PSmemory_2_0_arlock         (io_PSmemory_2_0_arlock),
      .io_PSmemory_2_0_arvalid        (io_PSmemory_2_0_arvalid),
      .io_PSmemory_2_0_arready        (io_PSmemory_2_0_arready),
      //.io_PSmemory_2_0_rid            (io_PSmemory_2_0_rid),
      .io_PSmemory_2_0_rdata          (io_PSmemory_2_0_rdata),
      .io_PSmemory_2_0_rresp          (io_PSmemory_2_0_rresp),
      .io_PSmemory_2_0_rlast          (io_PSmemory_2_0_rlast),
      .io_PSmemory_2_0_rvalid         (io_PSmemory_2_0_rvalid),
      .io_PSmemory_2_0_rready         (io_PSmemory_2_0_rready),
      
      //.io_PSmemory_2_1_awid           (io_PSmemory_2_1_awid),
      .io_PSmemory_2_1_awaddr         (io_PSmemory_2_1_awaddr),
      .io_PSmemory_2_1_awlen          (io_PSmemory_2_1_awlen),
      .io_PSmemory_2_1_awsize         (io_PSmemory_2_1_awsize),
      .io_PSmemory_2_1_awburst        (io_PSmemory_2_1_awburst),
      .io_PSmemory_2_1_awlock         (io_PSmemory_2_1_awlock),
      .io_PSmemory_2_1_awvalid        (io_PSmemory_2_1_awvalid),
      .io_PSmemory_2_1_awready        (io_PSmemory_2_1_awready),
      .io_PSmemory_2_1_wdata          (io_PSmemory_2_1_wdata),
      .io_PSmemory_2_1_wstrb          (io_PSmemory_2_1_wstrb),
      .io_PSmemory_2_1_wlast          (io_PSmemory_2_1_wlast),
      .io_PSmemory_2_1_wvalid         (io_PSmemory_2_1_wvalid),
      .io_PSmemory_2_1_wready         (io_PSmemory_2_1_wready),
      //.io_PSmemory_2_1_bid            (io_PSmemory_2_1_bid),
      .io_PSmemory_2_1_bresp          (io_PSmemory_2_1_bresp),
      .io_PSmemory_2_1_bvalid         (io_PSmemory_2_1_bvalid),
      .io_PSmemory_2_1_bready         (io_PSmemory_2_1_bready),
      //.io_PSmemory_2_1_arid           (io_PSmemory_2_1_arid),
      .io_PSmemory_2_1_araddr         (io_PSmemory_2_1_araddr),
      .io_PSmemory_2_1_arlen          (io_PSmemory_2_1_arlen),
      .io_PSmemory_2_1_arsize         (io_PSmemory_2_1_arsize),
      .io_PSmemory_2_1_arburst        (io_PSmemory_2_1_arburst),
      .io_PSmemory_2_1_arlock         (io_PSmemory_2_1_arlock),
      .io_PSmemory_2_1_arvalid        (io_PSmemory_2_1_arvalid),
      .io_PSmemory_2_1_arready        (io_PSmemory_2_1_arready),
      //.io_PSmemory_2_1_rid            (io_PSmemory_2_1_rid),
      .io_PSmemory_2_1_rdata          (io_PSmemory_2_1_rdata),
      .io_PSmemory_2_1_rresp          (io_PSmemory_2_1_rresp),
      .io_PSmemory_2_1_rlast          (io_PSmemory_2_1_rlast),
      .io_PSmemory_2_1_rvalid         (io_PSmemory_2_1_rvalid),
      .io_PSmemory_2_1_rready         (io_PSmemory_2_1_rready),
      
      //.io_PSmemory_3_0_awid           (io_PSmemory_3_0_awid),
      .io_PSmemory_3_0_awaddr         (io_PSmemory_3_0_awaddr),
      .io_PSmemory_3_0_awlen          (io_PSmemory_3_0_awlen),
      .io_PSmemory_3_0_awsize         (io_PSmemory_3_0_awsize),
      .io_PSmemory_3_0_awburst        (io_PSmemory_3_0_awburst),
      .io_PSmemory_3_0_awlock         (io_PSmemory_3_0_awlock),
      .io_PSmemory_3_0_awvalid        (io_PSmemory_3_0_awvalid),
      .io_PSmemory_3_0_awready        (io_PSmemory_3_0_awready),
      .io_PSmemory_3_0_wdata          (io_PSmemory_3_0_wdata),
      .io_PSmemory_3_0_wstrb          (io_PSmemory_3_0_wstrb),
      .io_PSmemory_3_0_wlast          (io_PSmemory_3_0_wlast),
      .io_PSmemory_3_0_wvalid         (io_PSmemory_3_0_wvalid),
      .io_PSmemory_3_0_wready         (io_PSmemory_3_0_wready),
      //.io_PSmemory_3_0_bid            (io_PSmemory_3_0_bid),
      .io_PSmemory_3_0_bresp          (io_PSmemory_3_0_bresp),
      .io_PSmemory_3_0_bvalid         (io_PSmemory_3_0_bvalid),
      .io_PSmemory_3_0_bready         (io_PSmemory_3_0_bready),
      //.io_PSmemory_3_0_arid           (io_PSmemory_3_0_arid),
      .io_PSmemory_3_0_araddr         (io_PSmemory_3_0_araddr),
      .io_PSmemory_3_0_arlen          (io_PSmemory_3_0_arlen),
      .io_PSmemory_3_0_arsize         (io_PSmemory_3_0_arsize),
      .io_PSmemory_3_0_arburst        (io_PSmemory_3_0_arburst),
      .io_PSmemory_3_0_arlock         (io_PSmemory_3_0_arlock),
      .io_PSmemory_3_0_arvalid        (io_PSmemory_3_0_arvalid),
      .io_PSmemory_3_0_arready        (io_PSmemory_3_0_arready),
      //.io_PSmemory_3_0_rid            (io_PSmemory_3_0_rid),
      .io_PSmemory_3_0_rdata          (io_PSmemory_3_0_rdata),
      .io_PSmemory_3_0_rresp          (io_PSmemory_3_0_rresp),
      .io_PSmemory_3_0_rlast          (io_PSmemory_3_0_rlast),
      .io_PSmemory_3_0_rvalid         (io_PSmemory_3_0_rvalid),
      .io_PSmemory_3_0_rready         (io_PSmemory_3_0_rready),
      
      //.io_PSmemory_3_1_awid           (io_PSmemory_3_1_awid),
      .io_PSmemory_3_1_awaddr         (io_PSmemory_3_1_awaddr),
      .io_PSmemory_3_1_awlen          (io_PSmemory_3_1_awlen),
      .io_PSmemory_3_1_awsize         (io_PSmemory_3_1_awsize),
      .io_PSmemory_3_1_awburst        (io_PSmemory_3_1_awburst),
      .io_PSmemory_3_1_awlock         (io_PSmemory_3_1_awlock),
      .io_PSmemory_3_1_awvalid        (io_PSmemory_3_1_awvalid),
      .io_PSmemory_3_1_awready        (io_PSmemory_3_1_awready),
      .io_PSmemory_3_1_wdata          (io_PSmemory_3_1_wdata),
      .io_PSmemory_3_1_wstrb          (io_PSmemory_3_1_wstrb),
      .io_PSmemory_3_1_wlast          (io_PSmemory_3_1_wlast),
      .io_PSmemory_3_1_wvalid         (io_PSmemory_3_1_wvalid),
      .io_PSmemory_3_1_wready         (io_PSmemory_3_1_wready),
      //.io_PSmemory_3_1_bid            (io_PSmemory_3_1_bid),
      .io_PSmemory_3_1_bresp          (io_PSmemory_3_1_bresp),
      .io_PSmemory_3_1_bvalid         (io_PSmemory_3_1_bvalid),
      .io_PSmemory_3_1_bready         (io_PSmemory_3_1_bready),
      //.io_PSmemory_3_1_arid           (io_PSmemory_3_1_arid),
      .io_PSmemory_3_1_araddr         (io_PSmemory_3_1_araddr),
      .io_PSmemory_3_1_arlen          (io_PSmemory_3_1_arlen),
      .io_PSmemory_3_1_arsize         (io_PSmemory_3_1_arsize),
      .io_PSmemory_3_1_arburst        (io_PSmemory_3_1_arburst),
      .io_PSmemory_3_1_arlock         (io_PSmemory_3_1_arlock),
      .io_PSmemory_3_1_arvalid        (io_PSmemory_3_1_arvalid),
      .io_PSmemory_3_1_arready        (io_PSmemory_3_1_arready),
      //.io_PSmemory_3_1_rid            (io_PSmemory_3_1_rid),
      .io_PSmemory_3_1_rdata          (io_PSmemory_3_1_rdata),
      .io_PSmemory_3_1_rresp          (io_PSmemory_3_1_rresp),
      .io_PSmemory_3_1_rlast          (io_PSmemory_3_1_rlast),
      .io_PSmemory_3_1_rvalid         (io_PSmemory_3_1_rvalid),
      .io_PSmemory_3_1_rready         (io_PSmemory_3_1_rready),
      
      .io_PSMemory_araddr         (io_PSmempory_ar_bits_araddr),
      .io_PSMemory_arburst        (io_PSmempory_ar_bits_arburst),
      .io_PSMemory_arcache        (),
      .io_PSMemory_arid           ({2'd0, io_PSmempory_ar_bits_arid}),
      .io_PSMemory_arlen          (io_PSmempory_ar_bits_arlen),
      .io_PSMemory_arlock         (io_PSmempory_ar_bits_arlock),
      .io_PSMemory_arprot         (),
      .io_PSMemory_arqos          (),
      .io_PSMemory_arready        (io_PSmempory_ar_ready),
      .io_PSMemory_arsize         (io_PSmempory_ar_bits_arsize),
      .io_PSMemory_arvalid        (io_PSmempory_ar_valid),
      .io_PSMemory_awaddr         (io_PSmempory_aw_bits_awaddr),
      .io_PSMemory_awburst        (io_PSmempory_aw_bits_awburst),
      .io_PSMemory_awcache        (),
      .io_PSMemory_awid           ({2'd0, io_PSmempory_aw_bits_awid}),
      .io_PSMemory_awlen          (io_PSmempory_aw_bits_awlen),
      .io_PSMemory_awlock         (io_PSmempory_aw_bits_awlock),
      .io_PSMemory_awprot         (),
      .io_PSMemory_awqos          (),
      .io_PSMemory_awready        (io_PSmempory_aw_ready),
      .io_PSMemory_awsize         (io_PSmempory_aw_bits_awsize),
      .io_PSMemory_awvalid        (io_PSmempory_aw_valid),
      .io_PSMemory_bid            (io_PSmempory_b_bits_bid),
      .io_PSMemory_bready         (io_PSmempory_b_ready),
      .io_PSMemory_bresp          (io_PSmempory_b_bits_bresp),
      .io_PSMemory_bvalid         (io_PSmempory_b_valid),
      .io_PSMemory_rdata          (io_PSmempory_r_bits_rdata),
      .io_PSMemory_rid            (io_PSmempory_r_bits_rid),
      .io_PSMemory_rlast          (io_PSmempory_r_bits_rlast),
      .io_PSMemory_rready         (io_PSmempory_r_ready),
      .io_PSMemory_rresp          (),
      .io_PSMemory_rvalid         (io_PSmempory_r_valid),
      .io_PSMemory_wdata          (io_PSmempory_w_bits_wdata),
      .io_PSMemory_wlast          (io_PSmempory_w_bits_wlast),
      .io_PSMemory_wready         (io_PSmempory_w_ready),
      .io_PSMemory_wstrb          (io_PSmempory_w_bits_wstrb),
      .io_PSMemory_wvalid         (io_PSmempory_w_valid),

      .io_PSMemory_1_araddr         (io_PSmempory_1_ar_bits_araddr),
      .io_PSMemory_1_arburst        (io_PSmempory_1_ar_bits_arburst),
      .io_PSMemory_1_arid           ({2'd1, io_PSmempory_1_ar_bits_arid}),
      .io_PSMemory_1_arlen          (io_PSmempory_1_ar_bits_arlen),
      .io_PSMemory_1_arlock         (io_PSmempory_1_ar_bits_arlock),
      .io_PSMemory_1_arready        (io_PSmempory_1_ar_ready),
      .io_PSMemory_1_arsize         (io_PSmempory_1_ar_bits_arsize),
      .io_PSMemory_1_arvalid        (io_PSmempory_1_ar_valid),
      .io_PSMemory_1_awaddr         (io_PSmempory_1_aw_bits_awaddr),
      .io_PSMemory_1_awburst        (io_PSmempory_1_aw_bits_awburst),
      .io_PSMemory_1_awid           ({2'd1, io_PSmempory_1_aw_bits_awid}),
      .io_PSMemory_1_awlen          (io_PSmempory_1_aw_bits_awlen),
      .io_PSMemory_1_awlock         (io_PSmempory_1_aw_bits_awlock),
      .io_PSMemory_1_awready        (io_PSmempory_1_aw_ready),
      .io_PSMemory_1_awsize         (io_PSmempory_1_aw_bits_awsize),
      .io_PSMemory_1_awvalid        (io_PSmempory_1_aw_valid),
      .io_PSMemory_1_bid            (io_PSmempory_1_b_bits_bid),
      .io_PSMemory_1_bready         (io_PSmempory_1_b_ready),
      .io_PSMemory_1_bresp          (io_PSmempory_1_b_bits_bresp),
      .io_PSMemory_1_bvalid         (io_PSmempory_1_b_valid),
      .io_PSMemory_1_rdata          (io_PSmempory_1_r_bits_rdata),
      .io_PSMemory_1_rid            (io_PSmempory_1_r_bits_rid),
      .io_PSMemory_1_rlast          (io_PSmempory_1_r_bits_rlast),
      .io_PSMemory_1_rready         (io_PSmempory_1_r_ready),
      .io_PSMemory_1_rvalid         (io_PSmempory_1_r_valid),
      .io_PSMemory_1_wdata          (io_PSmempory_1_w_bits_wdata),
      .io_PSMemory_1_wlast          (io_PSmempory_1_w_bits_wlast),
      .io_PSMemory_1_wready         (io_PSmempory_1_w_ready),
      .io_PSMemory_1_wstrb          (io_PSmempory_1_w_bits_wstrb),
      .io_PSMemory_1_wvalid         (io_PSmempory_1_w_valid),

      .io_PSMemory_2_araddr         (io_PSmempory_2_ar_bits_araddr),
      .io_PSMemory_2_arburst        (io_PSmempory_2_ar_bits_arburst),
      .io_PSMemory_2_arid           ({2'd2, io_PSmempory_2_ar_bits_arid}),
      .io_PSMemory_2_arlen          (io_PSmempory_2_ar_bits_arlen),
      .io_PSMemory_2_arlock         (io_PSmempory_2_ar_bits_arlock),
      .io_PSMemory_2_arready        (io_PSmempory_2_ar_ready),
      .io_PSMemory_2_arsize         (io_PSmempory_2_ar_bits_arsize),
      .io_PSMemory_2_arvalid        (io_PSmempory_2_ar_valid),
      .io_PSMemory_2_awaddr         (io_PSmempory_2_aw_bits_awaddr),
      .io_PSMemory_2_awburst        (io_PSmempory_2_aw_bits_awburst),
      .io_PSMemory_2_awid           ({2'd2, io_PSmempory_2_aw_bits_awid}),
      .io_PSMemory_2_awlen          (io_PSmempory_2_aw_bits_awlen),
      .io_PSMemory_2_awlock         (io_PSmempory_2_aw_bits_awlock),
      .io_PSMemory_2_awready        (io_PSmempory_2_aw_ready),
      .io_PSMemory_2_awsize         (io_PSmempory_2_aw_bits_awsize),
      .io_PSMemory_2_awvalid        (io_PSmempory_2_aw_valid),
      .io_PSMemory_2_bid            (io_PSmempory_2_b_bits_bid),
      .io_PSMemory_2_bready         (io_PSmempory_2_b_ready),
      .io_PSMemory_2_bresp          (io_PSmempory_2_b_bits_bresp),
      .io_PSMemory_2_bvalid         (io_PSmempory_2_b_valid),
      .io_PSMemory_2_rdata          (io_PSmempory_2_r_bits_rdata),
      .io_PSMemory_2_rid            (io_PSmempory_2_r_bits_rid),
      .io_PSMemory_2_rlast          (io_PSmempory_2_r_bits_rlast),
      .io_PSMemory_2_rready         (io_PSmempory_2_r_ready),
      .io_PSMemory_2_rvalid         (io_PSmempory_2_r_valid),
      .io_PSMemory_2_wdata          (io_PSmempory_2_w_bits_wdata),
      .io_PSMemory_2_wlast          (io_PSmempory_2_w_bits_wlast),
      .io_PSMemory_2_wready         (io_PSmempory_2_w_ready),
      .io_PSMemory_2_wstrb          (io_PSmempory_2_w_bits_wstrb),
      .io_PSMemory_2_wvalid         (io_PSmempory_2_w_valid),

      .io_PSMemory_3_araddr         (io_PSmempory_3_ar_bits_araddr),
      .io_PSMemory_3_arburst        (io_PSmempory_3_ar_bits_arburst),
      .io_PSMemory_3_arid           ({2'd3, io_PSmempory_3_ar_bits_arid}),
      .io_PSMemory_3_arlen          (io_PSmempory_3_ar_bits_arlen),
      .io_PSMemory_3_arlock         (io_PSmempory_3_ar_bits_arlock),
      .io_PSMemory_3_arready        (io_PSmempory_3_ar_ready),
      .io_PSMemory_3_arsize         (io_PSmempory_3_ar_bits_arsize),
      .io_PSMemory_3_arvalid        (io_PSmempory_3_ar_valid),
      .io_PSMemory_3_awaddr         (io_PSmempory_3_aw_bits_awaddr),
      .io_PSMemory_3_awburst        (io_PSmempory_3_aw_bits_awburst),
      .io_PSMemory_3_awid           ({2'd3, io_PSmempory_3_aw_bits_awid}),
      .io_PSMemory_3_awlen          (io_PSmempory_3_aw_bits_awlen),
      .io_PSMemory_3_awlock         (io_PSmempory_3_aw_bits_awlock),
      .io_PSMemory_3_awready        (io_PSmempory_3_aw_ready),
      .io_PSMemory_3_awsize         (io_PSmempory_3_aw_bits_awsize),
      .io_PSMemory_3_awvalid        (io_PSmempory_3_aw_valid),
      .io_PSMemory_3_bid            (io_PSmempory_3_b_bits_bid),
      .io_PSMemory_3_bready         (io_PSmempory_3_b_ready),
      .io_PSMemory_3_bresp          (io_PSmempory_3_b_bits_bresp),
      .io_PSMemory_3_bvalid         (io_PSmempory_3_b_valid),
      .io_PSMemory_3_rdata          (io_PSmempory_3_r_bits_rdata),
      .io_PSMemory_3_rid            (io_PSmempory_3_r_bits_rid),
      .io_PSMemory_3_rlast          (io_PSmempory_3_r_bits_rlast),
      .io_PSMemory_3_rready         (io_PSmempory_3_r_ready),
      .io_PSMemory_3_rvalid         (io_PSmempory_3_r_valid),
      .io_PSMemory_3_wdata          (io_PSmempory_3_w_bits_wdata),
      .io_PSMemory_3_wlast          (io_PSmempory_3_w_bits_wlast),
      .io_PSMemory_3_wready         (io_PSmempory_3_w_ready),
      .io_PSMemory_3_wstrb          (io_PSmempory_3_w_bits_wstrb),
      .io_PSMemory_3_wvalid         (io_PSmempory_3_w_valid),

      .io_Re_memory_out_araddr         (io_Re_memory_out_ar_bits_araddr),
      .io_Re_memory_out_arburst        (io_Re_memory_out_ar_bits_arburst),
      .io_Re_memory_out_arid           (io_Re_memory_out_ar_bits_arid),
      .io_Re_memory_out_arlen          (io_Re_memory_out_ar_bits_arlen),
      .io_Re_memory_out_arlock         (io_Re_memory_out_ar_bits_arlock),
      .io_Re_memory_out_arready        (io_Re_memory_out_ar_ready),
      .io_Re_memory_out_arsize         (io_Re_memory_out_ar_bits_arsize),
      .io_Re_memory_out_arvalid        (io_Re_memory_out_ar_valid),
      .io_Re_memory_out_awaddr         (io_Re_memory_out_aw_bits_awaddr),
      .io_Re_memory_out_awburst        (io_Re_memory_out_aw_bits_awburst),
      .io_Re_memory_out_awid           (io_Re_memory_out_aw_bits_awid),
      .io_Re_memory_out_awlen          (io_Re_memory_out_aw_bits_awlen),
      .io_Re_memory_out_awlock         (io_Re_memory_out_aw_bits_awlock),
      .io_Re_memory_out_awready        (io_Re_memory_out_aw_ready),
      .io_Re_memory_out_awsize         (io_Re_memory_out_aw_bits_awsize),
      .io_Re_memory_out_awvalid        (io_Re_memory_out_aw_valid),
      .io_Re_memory_out_bid            (io_Re_memory_out_b_bits_bid),
      .io_Re_memory_out_bready         (io_Re_memory_out_b_ready),
      .io_Re_memory_out_bresp          (io_Re_memory_out_b_bits_bresp),
      .io_Re_memory_out_bvalid         (io_Re_memory_out_b_valid),
      .io_Re_memory_out_rdata          (io_Re_memory_out_r_bits_rdata),
      .io_Re_memory_out_rid            (io_Re_memory_out_r_bits_rid),
      .io_Re_memory_out_rlast          (io_Re_memory_out_r_bits_rlast),
      .io_Re_memory_out_rready         (io_Re_memory_out_r_ready),
      .io_Re_memory_out_rvalid         (io_Re_memory_out_r_valid),
      .io_Re_memory_out_wdata          (io_Re_memory_out_w_bits_wdata),
      .io_Re_memory_out_wlast          (io_Re_memory_out_w_bits_wlast),
      .io_Re_memory_out_wready         (io_Re_memory_out_w_ready),
      .io_Re_memory_out_wstrb          (io_Re_memory_out_w_bits_wstrb),
      .io_Re_memory_out_wvalid         (io_Re_memory_out_w_valid),

      .io_Re_memory_in_araddr         (io_Re_memory_in_ar_bits_araddr),
      .io_Re_memory_in_arburst        (io_Re_memory_in_ar_bits_arburst),
      .io_Re_memory_in_arid           (io_Re_memory_in_ar_bits_arid),
      .io_Re_memory_in_arlen          (io_Re_memory_in_ar_bits_arlen),
      .io_Re_memory_in_arlock         (io_Re_memory_in_ar_bits_arlock),
      .io_Re_memory_in_arready        (io_Re_memory_in_ar_ready),
      .io_Re_memory_in_arsize         (io_Re_memory_in_ar_bits_arsize),
      .io_Re_memory_in_arvalid        (io_Re_memory_in_ar_valid),
      .io_Re_memory_in_awaddr         (io_Re_memory_in_aw_bits_awaddr),
      .io_Re_memory_in_awburst        (io_Re_memory_in_aw_bits_awburst),
      .io_Re_memory_in_awid           (io_Re_memory_in_aw_bits_awid),
      .io_Re_memory_in_awlen          (io_Re_memory_in_aw_bits_awlen),
      .io_Re_memory_in_awlock         (io_Re_memory_in_aw_bits_awlock),
      .io_Re_memory_in_awready        (io_Re_memory_in_aw_ready),
      .io_Re_memory_in_awsize         (io_Re_memory_in_aw_bits_awsize),
      .io_Re_memory_in_awvalid        (io_Re_memory_in_aw_valid),
      .io_Re_memory_in_bid            (io_Re_memory_in_b_bits_bid),
      .io_Re_memory_in_bready         (io_Re_memory_in_b_ready),
      .io_Re_memory_in_bresp          (io_Re_memory_in_b_bits_bresp),
      .io_Re_memory_in_bvalid         (io_Re_memory_in_b_valid),
      .io_Re_memory_in_rdata          (io_Re_memory_in_r_bits_rdata),
      .io_Re_memory_in_rid            (io_Re_memory_in_r_bits_rid),
      .io_Re_memory_in_rlast          (io_Re_memory_in_r_bits_rlast),
      .io_Re_memory_in_rready         (io_Re_memory_in_r_ready),
      .io_Re_memory_in_rvalid         (io_Re_memory_in_r_valid),
      .io_Re_memory_in_wdata          (io_Re_memory_in_w_bits_wdata),
      .io_Re_memory_in_wlast          (io_Re_memory_in_w_bits_wlast),
      .io_Re_memory_in_wready         (io_Re_memory_in_w_ready),
      .io_Re_memory_in_wstrb          (io_Re_memory_in_w_bits_wstrb),
      .io_Re_memory_in_wvalid         (io_Re_memory_in_w_valid),

      .io_config_in_awaddr     (io_config_awaddr),
      .io_config_in_awvalid    (io_config_awvalid),
      .io_config_in_awready    (io_config_awready),
      .io_config_in_awlen      ('d0),
      .io_config_in_awsize     ('d2),
      .io_config_in_araddr     (io_config_araddr),
      .io_config_in_arvalid    (io_config_arvalid),
      .io_config_in_arready    (io_config_arready),
      .io_config_in_wdata      (io_config_wdata),
      .io_config_in_wstrb      (io_config_wstrb),
      .io_config_in_wlast      (1'b1),
      .io_config_in_wvalid     (io_config_wvalid),
      .io_config_in_wready     (io_config_wready),
      .io_config_in_rdata      (io_config_rdata),
      .io_config_in_rresp      (io_config_rresp),
      .io_config_in_rvalid     (io_config_rvalid),
      .io_config_in_rready     (io_config_rready),
      .io_config_in_bresp      (io_config_bresp),
      .io_config_in_bvalid     (io_config_bvalid),
      .io_config_in_bready     (io_config_bready),

      .io_config_out_awaddr     (bfs_io_config_awaddr),
      .io_config_out_awvalid    (bfs_io_config_awvalid),
      .io_config_out_awready    (bfs_io_config_awready),
      .io_config_out_araddr     (bfs_io_config_araddr),
      .io_config_out_arvalid    (bfs_io_config_arvalid),
      .io_config_out_arready    (bfs_io_config_arready),
      .io_config_out_wdata      (bfs_io_config_wdata),
      .io_config_out_wstrb      (bfs_io_config_wstrb),
      .io_config_out_wvalid     (bfs_io_config_wvalid),
      .io_config_out_wready     (bfs_io_config_wready),
      .io_config_out_rdata      (bfs_io_config_rdata),
      .io_config_out_rresp      (bfs_io_config_rresp),
      .io_config_out_rvalid     (bfs_io_config_rvalid),
      .io_config_out_rready     (bfs_io_config_rready),
      .io_config_out_bresp      (bfs_io_config_bresp),
      .io_config_out_bvalid     (bfs_io_config_bvalid),
      .io_config_out_bready     (bfs_io_config_bready)
    );

    BFS_ps u_BFS(
      .clock                (gt_txusrclk),
      .reset                (peripheral_reset),
      .io_config_awaddr     (bfs_io_config_awaddr),
      .io_config_awvalid    (bfs_io_config_awvalid),
      .io_config_awready    (bfs_io_config_awready),
      .io_config_araddr     (bfs_io_config_araddr),
      .io_config_arvalid    (bfs_io_config_arvalid),
      .io_config_arready    (bfs_io_config_arready),
      .io_config_wdata      (bfs_io_config_wdata),
      .io_config_wstrb      (bfs_io_config_wstrb),
      .io_config_wvalid     (bfs_io_config_wvalid),
      .io_config_wready     (bfs_io_config_wready),
      .io_config_rdata      (bfs_io_config_rdata),
      .io_config_rresp      (bfs_io_config_rresp),
      .io_config_rvalid     (bfs_io_config_rvalid),
      .io_config_rready     (bfs_io_config_rready),
      .io_config_bresp      (bfs_io_config_bresp),
      .io_config_bvalid     (bfs_io_config_bvalid),
      .io_config_bready     (bfs_io_config_bready),
      .io_PLmemory_0_aw_bits_awaddr   (io_PLmemory_0_awaddr),
      .io_PLmemory_0_aw_bits_awid     (io_PLmemory_0_awid),
      .io_PLmemory_0_aw_bits_awlen    (io_PLmemory_0_awlen),
      .io_PLmemory_0_aw_bits_awsize   (io_PLmemory_0_awsize),
      .io_PLmemory_0_aw_bits_awburst  (io_PLmemory_0_awburst),
      .io_PLmemory_0_aw_bits_awlock   (io_PLmemory_0_awlock),
      .io_PLmemory_0_aw_valid  (io_PLmemory_0_awvalid),
      .io_PLmemory_0_aw_ready  (io_PLmemory_0_awready),
      .io_PLmemory_0_ar_bits_araddr   (io_PLmemory_0_araddr),
      .io_PLmemory_0_ar_bits_arid     (io_PLmemory_0_arid),
      .io_PLmemory_0_ar_bits_arlen    (io_PLmemory_0_arlen),
      .io_PLmemory_0_ar_bits_arsize   (io_PLmemory_0_arsize),
      .io_PLmemory_0_ar_bits_arburst  (io_PLmemory_0_arburst),
      .io_PLmemory_0_ar_bits_arlock   (io_PLmemory_0_arlock),
      .io_PLmemory_0_ar_valid  (io_PLmemory_0_arvalid),
      .io_PLmemory_0_ar_ready  (io_PLmemory_0_arready),
      .io_PLmemory_0_w_bits_wdata    (io_PLmemory_0_wdata),
      .io_PLmemory_0_w_bits_wstrb    (io_PLmemory_0_wstrb),
      .io_PLmemory_0_w_bits_wlast    (io_PLmemory_0_wlast),
      .io_PLmemory_0_w_valid   (io_PLmemory_0_wvalid),
      .io_PLmemory_0_w_ready   (io_PLmemory_0_wready),
      .io_PLmemory_0_r_bits_rdata    (io_PLmemory_0_rdata),
      .io_PLmemory_0_r_bits_rid      (io_PLmemory_0_rid),
      .io_PLmemory_0_r_bits_rlast    (io_PLmemory_0_rlast),
      //.io_PLmemory_0_r_bits_rresp    (io_PLmemory_0_rresp),
      .io_PLmemory_0_r_valid   (io_PLmemory_0_rvalid),
      .io_PLmemory_0_r_ready   (io_PLmemory_0_rready),
      .io_PLmemory_0_b_bits_bresp    (io_PLmemory_0_bresp),
      .io_PLmemory_0_b_bits_bid      (io_PLmemory_0_bid),
      .io_PLmemory_0_b_valid   (io_PLmemory_0_bvalid),
      .io_PLmemory_0_b_ready   (io_PLmemory_0_bready),
      .io_PLmemory_1_aw_bits_awaddr   (io_PLmemory_1_awaddr),
      .io_PLmemory_1_aw_bits_awid     (io_PLmemory_1_awid),
      .io_PLmemory_1_aw_bits_awlen    (io_PLmemory_1_awlen),
      .io_PLmemory_1_aw_bits_awsize   (io_PLmemory_1_awsize),
      .io_PLmemory_1_aw_bits_awburst  (io_PLmemory_1_awburst),
      .io_PLmemory_1_aw_bits_awlock   (io_PLmemory_1_awlock),
      .io_PLmemory_1_aw_valid  (io_PLmemory_1_awvalid),
      .io_PLmemory_1_aw_ready  (io_PLmemory_1_awready),
      .io_PLmemory_1_ar_bits_araddr   (io_PLmemory_1_araddr),
      .io_PLmemory_1_ar_bits_arid     (io_PLmemory_1_arid),
      .io_PLmemory_1_ar_bits_arlen    (io_PLmemory_1_arlen),
      .io_PLmemory_1_ar_bits_arsize   (io_PLmemory_1_arsize),
      .io_PLmemory_1_ar_bits_arburst  (io_PLmemory_1_arburst),
      .io_PLmemory_1_ar_bits_arlock   (io_PLmemory_1_arlock),
      .io_PLmemory_1_ar_valid  (io_PLmemory_1_arvalid),
      .io_PLmemory_1_ar_ready  (io_PLmemory_1_arready),
      .io_PLmemory_1_w_bits_wdata    (io_PLmemory_1_wdata),
      .io_PLmemory_1_w_bits_wstrb    (io_PLmemory_1_wstrb),
      .io_PLmemory_1_w_bits_wlast    (io_PLmemory_1_wlast),
      .io_PLmemory_1_w_valid   (io_PLmemory_1_wvalid),
      .io_PLmemory_1_w_ready   (io_PLmemory_1_wready),
      .io_PLmemory_1_r_bits_rdata    (io_PLmemory_1_rdata),
      .io_PLmemory_1_r_bits_rid      (io_PLmemory_1_rid),
      .io_PLmemory_1_r_bits_rlast    (io_PLmemory_1_rlast),
      //.io_PLmemory_1_r_bits_rresp    (io_PLmemory_1_rresp),
      .io_PLmemory_1_r_valid   (io_PLmemory_1_rvalid),
      .io_PLmemory_1_r_ready   (io_PLmemory_1_rready),
      .io_PLmemory_1_b_bits_bresp    (io_PLmemory_1_bresp),
      .io_PLmemory_1_b_bits_bid      (io_PLmemory_1_bid),
      .io_PLmemory_1_b_valid   (io_PLmemory_1_bvalid),
      .io_PLmemory_1_b_ready   (io_PLmemory_1_bready),

      .io_PSmemory_0_aw_ready          (io_PSmempory_aw_ready),
      .io_PSmemory_0_aw_valid          (io_PSmempory_aw_valid),
      .io_PSmemory_0_aw_bits_awaddr    (io_PSmempory_aw_bits_awaddr),
      .io_PSmemory_0_aw_bits_awid      (io_PSmempory_aw_bits_awid),
      .io_PSmemory_0_aw_bits_awlen     (io_PSmempory_aw_bits_awlen),
      .io_PSmemory_0_aw_bits_awsize    (io_PSmempory_aw_bits_awsize),
      .io_PSmemory_0_aw_bits_awburst   (io_PSmempory_aw_bits_awburst),
      .io_PSmemory_0_aw_bits_awlock    (io_PSmempory_aw_bits_awlock),
      .io_PSmemory_0_ar_ready          (io_PSmempory_ar_ready),
      .io_PSmemory_0_ar_valid          (io_PSmempory_ar_valid),
      .io_PSmemory_0_ar_bits_araddr    (io_PSmempory_ar_bits_araddr),
      .io_PSmemory_0_ar_bits_arid      (io_PSmempory_ar_bits_arid),
      .io_PSmemory_0_ar_bits_arlen     (io_PSmempory_ar_bits_arlen),
      .io_PSmemory_0_ar_bits_arsize    (io_PSmempory_ar_bits_arsize),
      .io_PSmemory_0_ar_bits_arburst   (io_PSmempory_ar_bits_arburst),
      .io_PSmemory_0_ar_bits_arlock    (io_PSmempory_ar_bits_arlock),
      .io_PSmemory_0_w_ready           (io_PSmempory_w_ready),
      .io_PSmemory_0_w_valid           (io_PSmempory_w_valid),
      .io_PSmemory_0_w_bits_wdata      (io_PSmempory_w_bits_wdata),
      .io_PSmemory_0_w_bits_wstrb      (io_PSmempory_w_bits_wstrb),
      .io_PSmemory_0_w_bits_wlast      (io_PSmempory_w_bits_wlast),
      .io_PSmemory_0_r_ready           (io_PSmempory_r_ready),
      .io_PSmemory_0_r_valid           (io_PSmempory_r_valid),
      .io_PSmemory_0_r_bits_rdata      (io_PSmempory_r_bits_rdata),
      .io_PSmemory_0_r_bits_rid        (io_PSmempory_r_bits_rid),
      .io_PSmemory_0_r_bits_rlast      (io_PSmempory_r_bits_rlast),
      .io_PSmemory_0_b_ready           (io_PSmempory_b_ready),
      .io_PSmemory_0_b_valid           (io_PSmempory_b_valid),
      .io_PSmemory_0_b_bits_bresp      (io_PSmempory_b_bits_bresp),
      .io_PSmemory_0_b_bits_bid        (io_PSmempory_b_bits_bid),

      .io_PSmemory_1_aw_ready          (io_PSmempory_1_aw_ready),
      .io_PSmemory_1_aw_valid          (io_PSmempory_1_aw_valid),
      .io_PSmemory_1_aw_bits_awaddr    (io_PSmempory_1_aw_bits_awaddr),
      .io_PSmemory_1_aw_bits_awid      (io_PSmempory_1_aw_bits_awid),
      .io_PSmemory_1_aw_bits_awlen     (io_PSmempory_1_aw_bits_awlen),
      .io_PSmemory_1_aw_bits_awsize    (io_PSmempory_1_aw_bits_awsize),
      .io_PSmemory_1_aw_bits_awburst   (io_PSmempory_1_aw_bits_awburst),
      .io_PSmemory_1_aw_bits_awlock    (io_PSmempory_1_aw_bits_awlock),
      .io_PSmemory_1_ar_ready          (io_PSmempory_1_ar_ready),
      .io_PSmemory_1_ar_valid          (io_PSmempory_1_ar_valid),
      .io_PSmemory_1_ar_bits_araddr    (io_PSmempory_1_ar_bits_araddr),
      .io_PSmemory_1_ar_bits_arid      (io_PSmempory_1_ar_bits_arid),
      .io_PSmemory_1_ar_bits_arlen     (io_PSmempory_1_ar_bits_arlen),
      .io_PSmemory_1_ar_bits_arsize    (io_PSmempory_1_ar_bits_arsize),
      .io_PSmemory_1_ar_bits_arburst   (io_PSmempory_1_ar_bits_arburst),
      .io_PSmemory_1_ar_bits_arlock    (io_PSmempory_1_ar_bits_arlock),
      .io_PSmemory_1_w_ready           (io_PSmempory_1_w_ready),
      .io_PSmemory_1_w_valid           (io_PSmempory_1_w_valid),
      .io_PSmemory_1_w_bits_wdata      (io_PSmempory_1_w_bits_wdata),
      .io_PSmemory_1_w_bits_wstrb      (io_PSmempory_1_w_bits_wstrb),
      .io_PSmemory_1_w_bits_wlast      (io_PSmempory_1_w_bits_wlast),
      .io_PSmemory_1_r_ready           (io_PSmempory_1_r_ready),
      .io_PSmemory_1_r_valid           (io_PSmempory_1_r_valid),
      .io_PSmemory_1_r_bits_rdata      (io_PSmempory_1_r_bits_rdata),
      .io_PSmemory_1_r_bits_rid        (io_PSmempory_1_r_bits_rid),
      .io_PSmemory_1_r_bits_rlast      (io_PSmempory_1_r_bits_rlast),
      .io_PSmemory_1_b_ready           (io_PSmempory_1_b_ready),
      .io_PSmemory_1_b_valid           (io_PSmempory_1_b_valid),
      .io_PSmemory_1_b_bits_bresp      (io_PSmempory_1_b_bits_bresp),
      .io_PSmemory_1_b_bits_bid        (io_PSmempory_1_b_bits_bid),

      .io_PSmemory_2_aw_ready          (io_PSmempory_2_aw_ready),
      .io_PSmemory_2_aw_valid          (io_PSmempory_2_aw_valid),
      .io_PSmemory_2_aw_bits_awaddr    (io_PSmempory_2_aw_bits_awaddr),
      .io_PSmemory_2_aw_bits_awid      (io_PSmempory_2_aw_bits_awid),
      .io_PSmemory_2_aw_bits_awlen     (io_PSmempory_2_aw_bits_awlen),
      .io_PSmemory_2_aw_bits_awsize    (io_PSmempory_2_aw_bits_awsize),
      .io_PSmemory_2_aw_bits_awburst   (io_PSmempory_2_aw_bits_awburst),
      .io_PSmemory_2_aw_bits_awlock    (io_PSmempory_2_aw_bits_awlock),
      .io_PSmemory_2_ar_ready          (io_PSmempory_2_ar_ready),
      .io_PSmemory_2_ar_valid          (io_PSmempory_2_ar_valid),
      .io_PSmemory_2_ar_bits_araddr    (io_PSmempory_2_ar_bits_araddr),
      .io_PSmemory_2_ar_bits_arid      (io_PSmempory_2_ar_bits_arid),
      .io_PSmemory_2_ar_bits_arlen     (io_PSmempory_2_ar_bits_arlen),
      .io_PSmemory_2_ar_bits_arsize    (io_PSmempory_2_ar_bits_arsize),
      .io_PSmemory_2_ar_bits_arburst   (io_PSmempory_2_ar_bits_arburst),
      .io_PSmemory_2_ar_bits_arlock    (io_PSmempory_2_ar_bits_arlock),
      .io_PSmemory_2_w_ready           (io_PSmempory_2_w_ready),
      .io_PSmemory_2_w_valid           (io_PSmempory_2_w_valid),
      .io_PSmemory_2_w_bits_wdata      (io_PSmempory_2_w_bits_wdata),
      .io_PSmemory_2_w_bits_wstrb      (io_PSmempory_2_w_bits_wstrb),
      .io_PSmemory_2_w_bits_wlast      (io_PSmempory_2_w_bits_wlast),
      .io_PSmemory_2_r_ready           (io_PSmempory_2_r_ready),
      .io_PSmemory_2_r_valid           (io_PSmempory_2_r_valid),
      .io_PSmemory_2_r_bits_rdata      (io_PSmempory_2_r_bits_rdata),
      .io_PSmemory_2_r_bits_rid        (io_PSmempory_2_r_bits_rid),
      .io_PSmemory_2_r_bits_rlast      (io_PSmempory_2_r_bits_rlast),
      .io_PSmemory_2_b_ready           (io_PSmempory_2_b_ready),
      .io_PSmemory_2_b_valid           (io_PSmempory_2_b_valid),
      .io_PSmemory_2_b_bits_bresp      (io_PSmempory_2_b_bits_bresp),
      .io_PSmemory_2_b_bits_bid        (io_PSmempory_2_b_bits_bid),

      .io_PSmemory_3_aw_ready          (io_PSmempory_3_aw_ready),
      .io_PSmemory_3_aw_valid          (io_PSmempory_3_aw_valid),
      .io_PSmemory_3_aw_bits_awaddr    (io_PSmempory_3_aw_bits_awaddr),
      .io_PSmemory_3_aw_bits_awid      (io_PSmempory_3_aw_bits_awid),
      .io_PSmemory_3_aw_bits_awlen     (io_PSmempory_3_aw_bits_awlen),
      .io_PSmemory_3_aw_bits_awsize    (io_PSmempory_3_aw_bits_awsize),
      .io_PSmemory_3_aw_bits_awburst   (io_PSmempory_3_aw_bits_awburst),
      .io_PSmemory_3_aw_bits_awlock    (io_PSmempory_3_aw_bits_awlock),
      .io_PSmemory_3_ar_ready          (io_PSmempory_3_ar_ready),
      .io_PSmemory_3_ar_valid          (io_PSmempory_3_ar_valid),
      .io_PSmemory_3_ar_bits_araddr    (io_PSmempory_3_ar_bits_araddr),
      .io_PSmemory_3_ar_bits_arid      (io_PSmempory_3_ar_bits_arid),
      .io_PSmemory_3_ar_bits_arlen     (io_PSmempory_3_ar_bits_arlen),
      .io_PSmemory_3_ar_bits_arsize    (io_PSmempory_3_ar_bits_arsize),
      .io_PSmemory_3_ar_bits_arburst   (io_PSmempory_3_ar_bits_arburst),
      .io_PSmemory_3_ar_bits_arlock    (io_PSmempory_3_ar_bits_arlock),
      .io_PSmemory_3_w_ready           (io_PSmempory_3_w_ready),
      .io_PSmemory_3_w_valid           (io_PSmempory_3_w_valid),
      .io_PSmemory_3_w_bits_wdata      (io_PSmempory_3_w_bits_wdata),
      .io_PSmemory_3_w_bits_wstrb      (io_PSmempory_3_w_bits_wstrb),
      .io_PSmemory_3_w_bits_wlast      (io_PSmempory_3_w_bits_wlast),
      .io_PSmemory_3_r_ready           (io_PSmempory_3_r_ready),
      .io_PSmemory_3_r_valid           (io_PSmempory_3_r_valid),
      .io_PSmemory_3_r_bits_rdata      (io_PSmempory_3_r_bits_rdata),
      .io_PSmemory_3_r_bits_rid        (io_PSmempory_3_r_bits_rid),
      .io_PSmemory_3_r_bits_rlast      (io_PSmempory_3_r_bits_rlast),
      .io_PSmemory_3_b_ready           (io_PSmempory_3_b_ready),
      .io_PSmemory_3_b_valid           (io_PSmempory_3_b_valid),
      .io_PSmemory_3_b_bits_bresp      (io_PSmempory_3_b_bits_bresp),
      .io_PSmemory_3_b_bits_bid        (io_PSmempory_3_b_bits_bid),

      .io_Re_memory_out_aw_ready           (io_Re_memory_out_aw_ready),
      .io_Re_memory_out_aw_valid           (io_Re_memory_out_aw_valid),
      .io_Re_memory_out_aw_bits_awaddr     (io_Re_memory_out_aw_bits_awaddr),
      .io_Re_memory_out_aw_bits_awid       (io_Re_memory_out_aw_bits_awid),
      .io_Re_memory_out_aw_bits_awlen      (io_Re_memory_out_aw_bits_awlen),
      .io_Re_memory_out_aw_bits_awsize     (io_Re_memory_out_aw_bits_awsize),
      .io_Re_memory_out_aw_bits_awburst    (io_Re_memory_out_aw_bits_awburst),
      .io_Re_memory_out_aw_bits_awlock     (io_Re_memory_out_aw_bits_awlock),
      .io_Re_memory_out_ar_ready           (io_Re_memory_out_ar_ready),
      .io_Re_memory_out_ar_valid           (io_Re_memory_out_ar_valid),
      .io_Re_memory_out_ar_bits_araddr     (io_Re_memory_out_ar_bits_araddr),
      .io_Re_memory_out_ar_bits_arid       (io_Re_memory_out_ar_bits_arid),
      .io_Re_memory_out_ar_bits_arlen      (io_Re_memory_out_ar_bits_arlen),
      .io_Re_memory_out_ar_bits_arsize     (io_Re_memory_out_ar_bits_arsize),
      .io_Re_memory_out_ar_bits_arburst    (io_Re_memory_out_ar_bits_arburst),
      .io_Re_memory_out_ar_bits_arlock     (io_Re_memory_out_ar_bits_arlock),
      .io_Re_memory_out_w_ready            (io_Re_memory_out_w_ready),
      .io_Re_memory_out_w_valid            (io_Re_memory_out_w_valid),
      .io_Re_memory_out_w_bits_wdata       (io_Re_memory_out_w_bits_wdata),
      .io_Re_memory_out_w_bits_wstrb       (io_Re_memory_out_w_bits_wstrb),
      .io_Re_memory_out_w_bits_wlast       (io_Re_memory_out_w_bits_wlast),
      .io_Re_memory_out_r_ready            (io_Re_memory_out_r_ready),
      .io_Re_memory_out_r_valid            (io_Re_memory_out_r_valid),
      .io_Re_memory_out_r_bits_rdata       (io_Re_memory_out_r_bits_rdata),
      .io_Re_memory_out_r_bits_rid         (io_Re_memory_out_r_bits_rid),
      .io_Re_memory_out_r_bits_rlast       (io_Re_memory_out_r_bits_rlast),
      .io_Re_memory_out_b_ready            (io_Re_memory_out_b_ready),
      .io_Re_memory_out_b_valid            (io_Re_memory_out_b_valid),
      .io_Re_memory_out_b_bits_bresp       (io_Re_memory_out_b_bits_bresp),
      .io_Re_memory_out_b_bits_bid         (io_Re_memory_out_b_bits_bid),

      .io_Re_memory_in_aw_ready            (io_Re_memory_in_aw_ready),
      .io_Re_memory_in_aw_valid            (io_Re_memory_in_aw_valid),
      .io_Re_memory_in_aw_bits_awaddr      (io_Re_memory_in_aw_bits_awaddr),
      .io_Re_memory_in_aw_bits_awid        (io_Re_memory_in_aw_bits_awid),
      .io_Re_memory_in_aw_bits_awlen       (io_Re_memory_in_aw_bits_awlen),
      .io_Re_memory_in_aw_bits_awsize      (io_Re_memory_in_aw_bits_awsize),
      .io_Re_memory_in_aw_bits_awburst     (io_Re_memory_in_aw_bits_awburst),
      .io_Re_memory_in_aw_bits_awlock      (io_Re_memory_in_aw_bits_awlock),
      .io_Re_memory_in_ar_ready            (io_Re_memory_in_ar_ready),
      .io_Re_memory_in_ar_valid            (io_Re_memory_in_ar_valid),
      .io_Re_memory_in_ar_bits_araddr      (io_Re_memory_in_ar_bits_araddr),
      .io_Re_memory_in_ar_bits_arid        (io_Re_memory_in_ar_bits_arid),
      .io_Re_memory_in_ar_bits_arlen       (io_Re_memory_in_ar_bits_arlen),
      .io_Re_memory_in_ar_bits_arsize      (io_Re_memory_in_ar_bits_arsize),
      .io_Re_memory_in_ar_bits_arburst     (io_Re_memory_in_ar_bits_arburst),
      .io_Re_memory_in_ar_bits_arlock      (io_Re_memory_in_ar_bits_arlock),
      .io_Re_memory_in_w_ready             (io_Re_memory_in_w_ready),
      .io_Re_memory_in_w_valid             (io_Re_memory_in_w_valid),
      .io_Re_memory_in_w_bits_wdata        (io_Re_memory_in_w_bits_wdata),
      .io_Re_memory_in_w_bits_wstrb        (io_Re_memory_in_w_bits_wstrb),
      .io_Re_memory_in_w_bits_wlast        (io_Re_memory_in_w_bits_wlast),
      .io_Re_memory_in_r_ready             (io_Re_memory_in_r_ready),
      .io_Re_memory_in_r_valid             (io_Re_memory_in_r_valid),
      .io_Re_memory_in_r_bits_rdata        (io_Re_memory_in_r_bits_rdata),
      .io_Re_memory_in_r_bits_rid          (io_Re_memory_in_r_bits_rid),
      .io_Re_memory_in_r_bits_rlast        (io_Re_memory_in_r_bits_rlast),
      .io_Re_memory_in_b_ready             (io_Re_memory_in_b_ready),
      .io_Re_memory_in_b_valid             (io_Re_memory_in_b_valid),
      .io_Re_memory_in_b_bits_bresp        (io_Re_memory_in_b_bits_bresp),
      .io_Re_memory_in_b_bits_bid          (io_Re_memory_in_b_bits_bid)
    );
endmodule
